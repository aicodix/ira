-- code table generated from table_vector.txt by generate_table_vector_vhd.cc
--
-- Copyright 2019 Ahmet Inan <inan@aicodix.de>

use work.ldpc_scalar.all;
use work.ldpc_vector.all;

package table_vector is
	function init_vector_parities return vector_parities;
	function init_vector_counts return vector_counts;
	function init_vector_offsets return vector_offsets;
	function init_vector_shifts return vector_shifts;
end package;

package body table_vector is
	function init_vector_parities return vector_parities is
	begin
		return 180;
	end function;

	function init_vector_counts return vector_counts is
	begin
		return (
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
		others => count_scalar'low);
	end function;

	function init_vector_offsets return vector_offsets is
	begin
		return (
23,26,34,38,48,64,192,206,356,386,395,425,562,566,
22,33,47,54,167,179,288,333,347,381,527,529,703,707,
21,32,46,53,166,178,291,332,346,380,526,528,702,706,
4,31,51,63,174,176,240,300,356,374,525,536,712,716,
2,23,47,49,73,117,196,297,321,371,419,477,653,657,
6,13,29,36,156,161,186,250,329,366,455,518,542,546,
12,20,28,32,35,69,192,194,201,372,495,536,548,552,
7,9,16,47,165,174,288,297,354,462,462,534,710,714,
40,57,58,101,115,173,284,295,300,451,475,512,651,655,
2,3,44,49,55,163,244,271,343,413,484,523,699,703,
13,21,29,32,33,70,193,195,202,373,492,537,549,553,
14,17,50,54,56,89,207,236,249,416,421,466,592,596,
0,1,46,51,53,161,246,269,341,415,486,521,697,701,
4,9,19,25,39,118,219,231,349,399,432,446,575,579,
10,12,15,70,114,156,250,278,354,411,430,516,606,610,
43,56,57,132,151,170,211,260,312,380,492,521,668,672,
5,6,14,98,99,168,219,255,348,375,471,528,704,708,
7,19,48,53,79,141,259,309,351,384,439,508,615,619,
29,40,59,84,135,154,258,334,354,501,514,521,690,694,
6,10,17,45,65,86,226,266,328,415,440,446,622,626,
0,11,48,51,54,127,209,228,307,363,408,418,584,588,
14,24,25,39,64,143,244,339,340,365,424,458,600,604,
28,43,58,87,134,153,257,333,353,500,513,520,689,693,
16,32,33,40,48,86,212,221,357,385,392,466,568,572,
7,8,18,24,38,117,218,230,348,398,435,445,574,578,
3,17,29,54,127,176,236,287,307,396,487,537,663,667,
10,31,48,136,138,149,233,245,316,422,437,496,672,676,
4,7,12,96,97,170,217,253,350,373,469,530,706,710,
11,16,43,45,117,147,180,184,196,376,400,431,552,556,
6,8,9,30,122,161,188,204,341,363,368,456,544,548,
31,38,53,58,79,132,191,211,264,391,433,492,567,571,
2,23,24,94,94,146,223,259,274,427,438,454,630,634,
4,5,13,97,98,171,218,254,351,374,470,531,707,711,
1,9,14,26,41,124,181,238,278,361,376,507,541,716,
6,7,15,96,99,169,216,252,349,372,468,529,705,709,
5,8,11,29,121,160,191,207,340,362,371,459,547,551,
12,19,48,52,58,91,205,238,251,418,423,464,594,598,
23,33,42,80,110,153,187,260,297,440,454,531,616,620,
9,18,41,47,119,145,182,186,198,378,402,429,554,558,
1,39,46,98,111,152,278,312,321,458,499,535,634,638,
4,11,13,32,69,129,183,281,309,477,489,509,665,669,
23,34,44,55,164,176,289,334,344,382,524,530,700,704,
1,2,47,48,54,162,247,270,342,412,487,522,698,702,
3,31,57,59,101,106,233,269,286,466,482,513,642,646,
0,10,19,35,38,88,268,325,338,392,448,481,624,628,
18,30,43,61,72,105,241,275,344,410,421,501,597,601,
12,22,26,54,112,146,267,318,326,470,496,506,682,686,
21,35,40,82,108,155,185,262,299,442,452,529,618,622,
3,20,25,95,95,147,220,256,275,424,439,455,631,635,
1,19,31,52,125,178,238,285,305,398,485,539,661,665,
12,26,27,41,83,122,261,283,302,367,482,507,658,662,
22,25,33,37,51,67,195,205,359,385,394,424,561,565,
5,17,50,55,77,143,257,311,349,386,437,510,613,617,
20,35,45,52,165,177,290,335,345,383,525,531,701,705,
28,39,54,59,76,133,188,208,265,388,434,493,564,568,
14,24,25,43,81,120,263,281,300,365,480,505,656,660,
5,10,16,26,36,119,216,228,350,396,433,447,572,576,
4,15,31,38,158,163,184,248,331,364,453,516,540,544,
20,22,23,37,121,129,202,294,309,379,382,526,558,562,
21,24,32,36,50,66,194,204,358,384,393,427,560,564,
4,8,19,47,67,84,224,264,330,413,442,444,620,624,
16,28,41,63,74,107,243,273,346,408,423,503,599,603,
3,11,12,24,43,126,183,236,276,363,378,505,543,718,
18,34,35,42,50,84,214,223,359,387,394,464,570,574,
19,31,40,62,73,106,242,272,345,411,422,502,598,602,
3,21,33,45,63,93,225,227,229,388,405,489,581,585,
30,37,52,57,78,135,190,210,267,390,432,495,566,570,
1,22,46,48,72,116,199,296,320,370,418,476,652,656,
20,27,35,39,49,65,193,207,357,387,392,426,563,567,
29,36,55,56,77,134,189,209,266,389,435,494,565,569,
24,26,31,46,57,74,202,241,254,434,478,487,610,614,
7,30,50,62,173,179,243,303,359,373,524,539,715,719,
6,18,39,42,49,55,222,255,314,397,402,402,578,582,
19,32,35,43,51,85,215,220,356,384,395,465,571,575,
4,10,11,28,120,163,190,206,343,361,370,458,546,550,
7,14,30,37,157,162,187,251,330,367,452,519,543,547,
6,38,50,53,58,149,218,307,329,406,509,535,685,689,
3,28,43,79,129,158,199,335,338,405,445,518,694,698,
2,20,32,44,62,92,224,226,228,391,404,488,580,584,
8,17,40,46,118,144,181,185,197,377,401,428,553,557,
4,16,49,54,76,142,256,310,348,385,436,509,612,616,
3,37,44,96,109,154,276,314,323,456,497,533,632,636,
25,27,30,45,56,73,201,240,253,433,477,486,609,613,
6,29,49,61,172,178,242,302,358,372,527,538,714,718,
11,12,13,71,115,157,251,279,355,408,431,517,607,611,
7,19,36,43,50,52,223,252,315,398,403,403,579,583,
0,29,40,76,130,159,196,332,339,406,446,519,695,699,
15,23,31,34,35,68,193,195,200,375,494,539,551,555,
13,16,49,53,59,88,206,239,248,419,420,465,595,599,
2,8,17,33,36,90,270,327,336,394,450,483,626,630,
14,23,46,57,107,142,215,322,345,451,488,502,678,682,
20,21,22,39,123,131,200,292,311,377,380,524,556,560,
4,16,37,40,51,53,220,253,312,399,400,400,576,580,
2,9,49,50,52,125,211,230,305,361,410,416,586,590,
10,19,42,44,116,146,183,187,199,379,403,430,555,559,
15,20,47,58,104,143,212,323,346,448,489,503,679,683,
4,36,48,55,56,151,216,305,331,404,511,533,687,691,
5,37,49,52,57,148,217,306,328,405,508,534,684,688,
20,34,43,81,111,154,184,261,298,441,455,528,617,621,
9,14,15,69,113,159,249,277,353,410,429,519,605,609,
7,10,12,35,68,128,182,280,308,476,488,508,664,668,
16,41,44,52,54,165,214,234,275,414,431,442,590,594,
17,42,45,53,55,166,215,235,272,415,428,443,591,595,
7,11,18,46,66,87,227,267,329,412,441,447,623,627,
14,22,30,33,34,71,192,194,203,374,493,538,550,554,
25,35,37,81,110,138,188,290,293,391,470,472,646,650,
5,12,28,39,159,160,185,249,328,365,454,517,541,545,
20,21,23,38,122,130,203,295,310,376,383,527,559,563,
0,18,30,55,124,177,237,284,304,397,484,538,660,664,
15,25,26,36,65,140,245,336,341,366,425,459,601,605,
8,13,14,68,112,158,248,276,352,409,428,518,604,608,
5,17,38,41,48,54,221,254,313,396,401,401,577,581,
15,25,26,40,82,121,260,282,301,366,481,506,657,661,
8,29,50,136,138,151,235,247,318,420,439,498,674,678,
22,32,41,83,109,152,186,263,296,443,453,530,619,623,
11,28,49,137,139,150,234,246,317,423,438,497,673,677,
3,10,50,51,53,126,208,231,306,362,411,417,587,591,
1,29,57,59,103,104,235,271,284,464,480,515,640,644,
0,22,34,46,60,94,224,226,230,389,406,490,582,586,
6,18,51,52,78,140,258,308,350,387,438,511,614,618,
35,39,45,91,101,170,281,317,327,371,461,473,637,641,
17,33,34,41,49,87,213,222,358,386,393,467,569,573,
3,20,44,50,74,118,197,298,322,368,416,478,654,658,
25,27,28,47,58,75,203,242,255,435,479,484,611,615,
15,18,51,55,57,90,204,237,250,417,422,467,593,597,
12,21,44,59,105,140,213,320,347,449,490,500,676,680,
6,11,17,27,37,116,217,229,351,397,434,444,573,577,
7,9,10,31,123,162,189,205,342,360,369,457,545,549,
5,28,48,60,175,177,241,301,357,375,526,537,713,717,
19,40,47,53,55,164,213,233,274,413,430,441,589,593,
13,24,27,42,80,123,262,280,303,364,483,504,659,663,
4,10,17,44,166,175,289,298,355,463,463,535,711,715,
1,30,41,77,131,156,197,333,336,407,447,516,692,696,
2,16,28,53,126,179,239,286,306,399,486,536,662,666,
5,11,18,45,167,172,290,299,352,460,460,532,708,712,
13,23,27,55,113,147,264,319,327,471,497,507,683,687,
24,34,36,80,109,137,191,289,292,390,469,475,645,649,
0,38,45,97,110,155,277,315,320,457,498,534,633,637,
17,29,42,60,75,104,240,274,347,409,420,500,596,600,
1,23,35,47,61,95,225,227,231,390,407,491,583,587,
2,30,56,58,100,105,232,268,285,465,481,512,641,645,
24,26,29,44,59,72,200,243,252,432,476,485,608,612,
27,33,39,83,108,136,190,288,295,389,468,474,644,648,
31,42,57,86,133,152,256,332,352,503,512,523,688,692,
9,30,51,137,139,148,232,244,319,421,436,499,675,679,
1,11,16,32,39,89,269,326,339,393,449,482,625,629,
0,28,56,58,102,107,234,270,287,467,483,514,643,647,
2,36,47,99,108,153,279,313,322,459,496,532,635,639,
3,9,18,34,37,91,271,324,337,395,451,480,627,631,
0,8,13,25,40,127,180,237,277,360,379,506,540,719,
41,58,59,102,112,174,285,292,301,448,472,513,648,652,
43,56,57,100,114,172,287,294,303,450,474,515,650,654,
5,8,14,33,70,130,180,282,310,478,490,510,666,670,
1,22,27,93,93,145,222,258,273,426,437,453,629,633,
0,21,26,92,92,144,221,257,272,425,436,452,628,632,
34,38,44,90,100,169,280,316,326,370,460,472,636,640,
1,8,48,49,55,124,210,229,304,360,409,419,585,589,
2,10,15,27,42,125,182,239,279,362,377,504,542,717,
26,32,38,82,111,139,189,291,294,388,471,473,647,651,
18,43,46,52,54,167,212,232,273,412,429,440,588,592,
42,56,59,135,150,169,210,263,315,383,495,520,671,675,
0,21,45,51,75,119,198,299,323,369,417,479,655,659,
6,8,19,46,164,173,291,296,353,461,461,533,709,713,
5,9,16,44,64,85,225,265,331,414,443,445,621,625,
42,56,59,103,113,175,286,293,302,449,473,514,649,653,
12,26,27,37,66,141,246,337,342,367,426,456,602,606,
32,36,46,88,102,171,282,318,324,368,462,474,638,642,
6,9,15,34,71,131,181,283,311,479,491,511,667,671,
0,3,45,50,52,160,245,268,340,414,485,520,696,700,
30,41,56,85,132,155,259,335,355,502,515,522,691,695,
21,22,23,36,120,128,201,293,308,378,381,525,557,561,
13,24,27,38,67,142,247,338,343,364,427,457,603,607,
33,37,47,89,103,168,283,319,325,369,463,475,639,643,
40,57,58,133,148,171,208,261,313,381,493,522,669,673,
7,39,51,54,59,150,219,304,330,407,510,532,686,690,
2,31,42,78,128,157,198,334,337,404,444,517,693,697,
13,22,45,56,106,141,214,321,344,450,491,501,677,681,
14,20,24,52,114,144,265,316,324,468,498,504,680,684,
41,58,59,134,149,168,209,262,314,382,494,523,670,674,
15,21,25,53,115,145,266,317,325,469,499,505,681,685,
		others => 0);
	end function;

	function init_vector_shifts return vector_shifts is
	begin
		return (
11,0,39,87,42,16,73,0,56,0,63,75,0,0,
38,44,46,86,0,25,23,29,0,58,0,46,0,0,
38,44,46,86,0,25,22,29,0,58,0,46,0,0,
50,86,61,72,46,0,48,37,0,80,56,0,0,0,
76,58,89,82,79,0,82,0,74,18,47,0,0,0,
0,70,88,79,11,45,0,23,38,0,7,45,0,0,
0,55,68,87,12,17,0,24,51,0,48,74,0,0,
75,81,79,48,65,0,26,12,0,7,41,0,0,0,
51,42,3,51,0,43,67,0,18,43,0,13,0,0,
55,28,32,51,69,0,56,68,0,76,11,0,0,0,
0,55,68,13,87,17,0,24,51,0,49,74,0,0,
24,36,1,16,0,75,0,0,82,0,56,42,0,0,
55,28,31,50,69,0,55,68,0,75,10,0,0,0,
14,55,30,68,0,19,0,87,84,0,23,68,0,0,
6,11,16,0,42,48,0,7,77,27,0,34,0,0,
33,28,6,0,78,55,22,83,0,39,0,63,0,0,
88,85,41,11,73,0,19,39,0,44,62,0,0,0,
27,9,79,4,0,7,0,5,46,77,0,39,0,0,
20,88,14,56,29,0,74,0,42,28,0,24,0,0,
79,55,48,29,52,0,45,0,64,7,66,0,0,0,
72,45,0,62,75,12,6,0,36,70,0,46,0,0,
49,41,64,35,0,60,0,42,43,68,0,50,0,0,
20,87,14,55,29,0,74,0,42,28,0,24,0,0,
81,0,70,34,8,65,0,80,47,47,0,53,0,0,
13,55,30,68,0,19,0,87,84,0,22,68,0,0,
9,6,66,67,0,76,83,20,0,33,0,10,0,0,
15,48,2,0,76,84,67,27,0,17,58,0,0,0,
86,88,42,12,74,0,20,40,0,45,63,0,0,0,
9,0,50,3,42,79,83,20,0,0,85,42,0,0,
52,0,22,5,72,3,0,46,8,50,0,7,0,0,
0,20,53,45,50,12,75,0,69,0,41,16,0,0,
61,49,47,0,40,84,4,43,0,68,21,0,0,0,
89,86,42,12,74,0,20,40,0,45,63,0,0,0,
0,13,51,36,41,66,0,43,75,0,47,19,0,0,
88,85,41,74,11,0,20,40,0,45,63,0,0,0,
53,23,0,6,73,4,0,46,9,51,0,7,0,0,
25,36,2,17,0,75,1,0,82,0,56,43,0,0,
12,85,28,0,48,56,34,0,64,0,80,9,0,0,
10,0,51,3,42,80,83,20,0,0,85,43,0,0,
16,71,8,0,9,37,0,42,4,0,17,28,0,0,
27,46,69,71,16,0,84,55,0,53,0,52,0,0,
37,43,46,85,0,25,22,28,0,57,0,45,0,0,
55,28,31,51,69,0,55,68,0,76,10,0,0,0,
46,22,54,73,50,0,51,69,0,0,28,5,0,0,
75,14,26,56,49,0,0,44,74,3,0,24,0,0,
83,23,53,0,10,56,0,57,5,70,0,76,0,0,
47,2,5,44,77,0,13,49,0,88,10,0,0,0,
13,85,29,0,49,56,35,0,64,0,81,10,0,0,
61,50,47,0,40,84,5,44,0,69,21,0,0,0,
9,5,65,67,0,75,82,20,0,32,0,9,0,0,
82,57,71,49,68,0,12,59,0,13,0,54,0,0,
11,0,39,87,41,15,72,0,55,0,63,75,0,0,
27,9,78,3,0,6,0,4,46,76,0,38,0,0,
38,43,46,86,0,25,22,28,0,57,0,45,0,0,
0,19,52,44,50,11,75,0,68,0,40,15,0,0,
81,57,71,48,68,0,11,59,0,13,0,54,0,0,
13,54,30,67,0,18,0,87,83,0,22,67,0,0,
0,69,87,78,10,44,0,23,37,0,7,45,0,0,
21,0,82,50,71,14,0,1,23,82,0,6,0,0,
11,0,39,87,41,15,72,0,55,0,63,74,0,0,
79,55,47,28,51,0,45,0,63,7,65,0,0,0,
84,24,54,0,10,56,0,58,5,71,0,76,0,0,
0,13,52,37,41,66,0,44,76,0,47,20,0,0,
81,0,70,34,8,66,0,80,47,47,0,54,0,0,
83,23,54,0,10,56,0,58,5,70,0,76,0,0,
85,60,58,0,23,48,0,80,21,76,0,22,0,0,
0,20,53,45,50,11,75,0,68,0,41,15,0,0,
76,58,89,82,79,0,81,0,74,18,47,0,0,0,
12,0,39,87,42,16,73,0,56,0,64,75,0,0,
0,20,52,45,50,11,75,0,68,0,40,15,0,0,
33,33,39,30,10,0,12,36,0,0,13,26,0,0,
50,87,62,73,47,0,48,37,0,81,57,0,0,0,
5,63,53,0,70,87,0,45,4,24,0,80,0,0,
81,71,0,34,8,66,0,81,48,48,0,54,0,0,
53,0,22,6,73,3,0,46,8,51,0,7,0,0,
0,70,88,79,11,45,0,23,38,0,8,45,0,0,
19,72,75,46,63,0,7,12,0,27,0,61,0,0,
49,79,17,66,57,0,88,63,0,39,83,0,0,0,
85,60,58,0,23,48,0,80,21,75,0,22,0,0,
10,0,51,3,42,80,83,20,0,0,85,43,0,0,
27,9,78,3,0,6,0,4,46,76,0,38,0,0,
15,71,8,0,9,36,0,41,3,0,17,28,0,0,
33,32,39,30,10,0,12,36,0,0,13,26,0,0,
50,87,62,73,47,0,48,37,0,81,56,0,0,0,
6,17,11,0,42,48,0,7,77,28,0,34,0,0,
5,63,54,0,70,88,0,46,4,24,0,80,0,0,
50,79,18,67,57,0,89,64,0,39,83,0,0,0,
0,55,68,13,87,18,25,0,52,0,49,74,0,0,
25,37,2,17,0,76,1,0,83,0,57,43,0,0,
75,15,27,57,50,0,0,44,75,3,0,24,0,0,
58,81,89,19,14,0,54,0,47,13,1,0,0,0,
0,82,20,49,70,13,0,1,22,82,0,6,0,0,
5,63,53,0,69,87,0,45,4,23,0,80,0,0,
72,46,63,0,76,13,6,0,37,71,0,47,0,0,
10,0,51,4,43,80,83,20,0,0,85,43,0,0,
58,82,89,19,15,0,55,0,47,14,1,0,0,0,
20,73,76,46,64,0,8,13,0,28,0,62,0,0,
19,72,75,46,63,0,7,12,0,27,0,61,0,0,
13,85,28,0,48,56,35,0,64,0,80,10,0,0,
6,16,10,0,42,47,0,7,77,27,0,33,0,0,
26,46,69,70,16,0,84,55,0,53,0,52,0,0,
39,39,80,41,0,28,62,0,80,0,64,20,0,0,
39,39,80,41,0,28,62,0,81,0,65,20,0,0,
79,55,48,29,52,0,45,0,64,8,66,0,0,0,
0,55,68,13,87,17,25,0,51,0,49,74,0,0,
46,11,63,72,0,17,45,0,48,46,0,89,0,0,
0,70,88,78,10,45,0,23,38,0,7,45,0,0,
83,21,0,50,71,14,0,1,23,83,0,6,0,0,
9,5,65,66,0,75,82,20,0,32,0,9,0,0,
49,41,64,36,0,61,0,43,43,68,0,50,0,0,
6,16,10,0,42,47,0,7,77,27,0,33,0,0,
5,63,53,0,70,87,0,45,4,24,0,80,0,0,
81,57,71,49,68,0,12,59,0,13,0,54,0,0,
16,49,2,77,0,84,67,27,0,18,58,0,0,0,
13,86,29,0,49,57,35,0,65,0,81,10,0,0,
15,49,2,0,76,84,67,27,0,17,58,0,0,0,
72,46,63,0,76,13,7,0,37,71,0,47,0,0,
46,22,73,53,49,0,50,68,0,0,28,4,0,0,
86,60,58,0,24,48,81,0,21,76,0,22,0,0,
27,9,78,4,0,7,0,5,46,76,0,38,0,0,
55,63,26,12,0,14,0,5,73,47,0,19,0,0,
81,0,70,34,8,65,0,80,47,47,0,53,0,0,
76,59,0,82,79,0,82,0,74,19,48,0,0,0,
33,33,40,30,10,0,12,36,0,0,13,27,0,0,
24,36,1,16,0,75,1,0,82,0,56,42,0,0,
58,81,89,18,14,0,54,0,46,13,0,0,0,0,
13,54,30,67,0,19,0,87,83,0,22,68,0,0,
52,0,22,5,72,3,0,46,8,51,0,7,0,0,
50,87,62,73,46,0,48,37,0,80,56,0,0,0,
38,39,79,0,40,28,62,0,80,0,64,20,0,0,
82,72,57,49,69,0,12,60,0,14,0,55,0,0,
76,81,79,49,65,0,26,12,0,7,41,0,0,0,
49,78,17,66,56,0,88,63,0,38,82,0,0,0,
9,6,66,67,0,75,82,20,0,32,0,10,0,0,
75,80,78,48,64,0,25,11,0,7,41,0,0,0,
47,2,5,44,77,0,14,49,0,88,10,0,0,0,
46,11,63,72,0,17,44,0,48,46,0,88,0,0,
16,71,8,0,9,36,0,41,4,0,17,28,0,0,
83,23,53,0,9,56,0,57,4,70,0,76,0,0,
86,60,58,0,24,48,81,0,21,76,0,22,0,0,
46,22,54,73,50,0,51,69,0,0,28,5,0,0,
33,32,39,30,9,0,12,35,0,0,13,26,0,0,
45,11,62,71,0,17,44,0,47,46,0,88,0,0,
19,87,14,55,29,0,74,0,42,27,0,23,0,0,
16,49,2,77,0,85,68,28,0,18,59,0,0,0,
75,14,27,57,49,0,0,44,74,3,0,24,0,0,
47,23,74,54,50,0,51,69,0,0,28,5,0,0,
16,72,8,0,10,37,0,42,4,0,18,29,0,0,
75,15,27,57,50,0,0,45,75,3,0,25,0,0,
0,13,51,36,41,65,0,43,75,0,46,19,0,89,
50,41,2,50,0,42,66,0,17,43,0,12,0,0,
50,42,3,51,0,43,66,0,17,43,0,12,0,0,
27,47,69,71,16,0,85,55,0,53,0,52,0,0,
61,49,46,0,40,84,4,43,0,68,21,0,0,0,
61,49,46,0,40,84,4,43,0,68,21,0,0,0,
55,63,26,12,0,14,0,5,73,47,0,19,0,0,
72,46,63,0,75,13,6,0,37,71,0,46,0,0,
0,13,51,36,41,66,0,43,75,0,47,20,0,0,
46,12,63,72,0,17,45,0,48,47,0,89,0,0,
38,38,79,0,40,27,62,0,80,0,64,20,0,0,
34,7,28,0,79,56,23,83,0,39,0,64,0,0,
77,59,0,82,79,0,82,0,74,19,48,0,0,0,
75,81,78,48,65,0,25,12,0,7,41,0,0,0,
79,55,48,29,52,0,45,0,63,7,65,0,0,0,
50,3,41,50,0,42,66,0,17,43,0,12,0,0,
50,41,64,36,0,61,0,43,43,68,0,51,0,0,
56,64,26,13,0,14,0,5,74,48,0,19,0,0,
27,47,69,71,16,0,85,55,0,53,0,52,0,0,
28,54,31,50,69,0,55,68,0,75,10,0,0,0,
20,88,15,56,30,0,74,0,42,28,0,24,0,0,
0,82,20,50,71,14,0,1,23,82,0,6,0,0,
50,65,41,36,0,61,0,43,43,69,0,51,0,0,
56,64,26,13,0,15,0,5,74,48,0,19,0,0,
34,28,6,0,79,55,23,83,0,39,0,63,0,0,
19,72,75,46,63,0,7,13,0,27,0,62,0,0,
49,78,17,66,57,0,88,63,0,39,83,0,0,0,
58,81,89,19,14,0,54,0,47,13,0,0,0,0,
46,2,5,44,76,0,13,49,0,88,9,0,0,0,
34,28,6,0,79,56,23,83,0,39,0,63,0,0,
46,2,5,44,76,0,13,49,0,88,9,0,0,0,
		others => 0);
	end function;
end package body;
