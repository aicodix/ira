-- code table generated from table_vector.txt by generate_table_vector_vhd.cc
--
-- Copyright 2019 Ahmet Inan <inan@aicodix.de>

use work.ldpc_scalar.all;
use work.ldpc_vector.all;

package table_vector is
	function init_vector_parities return vector_parities;
	function init_vector_counts return vector_counts;
	function init_vector_offsets return vector_offsets;
	function init_vector_shifts return vector_shifts;
end package;

package body table_vector is
	function init_vector_parities return vector_parities is
	begin
		return 1080;
	end function;

	function init_vector_counts return vector_counts is
	begin
		return (
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
		others => count_scalar'low);
	end function;

	function init_vector_offsets return vector_offsets is
	begin
		return (
122,132,139,225,741,777,1202,1758,1869,2275,2282,3146,3338,3362,
26,114,219,246,309,331,1326,1531,1894,2381,2406,2414,3462,3486,
4,50,99,195,238,544,1624,1945,2018,2356,2704,2897,3760,3784,
123,130,140,233,725,785,1210,1766,1853,2259,2290,3154,3346,3370,
10,49,298,309,312,757,1259,1378,1837,2165,2458,2500,3514,3538,
125,196,278,317,1006,1058,1743,2008,2086,2292,3166,3180,4222,4246,
0,168,342,348,614,631,1410,1626,1711,2791,2903,3074,3847,3871,
124,131,141,234,726,786,1211,1767,1854,2260,2291,3155,3347,3371,
162,192,230,482,651,839,1141,1731,1754,2348,2811,2853,3867,3891,
137,211,248,494,664,935,1113,1574,1783,2654,2712,3173,3710,3734,
183,238,321,338,479,804,1131,1263,1584,2343,2601,2956,3399,3423,
0,52,85,145,260,767,1080,1421,1669,2160,2275,3030,3240,4319,
113,185,258,380,443,628,1460,1642,2079,2461,2540,3012,3596,3620,
135,209,246,492,662,933,1111,1572,1781,2652,2734,3171,3708,3732,
182,261,352,517,796,919,1551,1999,2119,3022,3079,3126,4135,4159,
5,16,282,311,313,973,1482,1629,2053,2475,2910,3133,4189,4213,
83,128,279,358,628,859,1292,1939,2078,2688,2949,3019,4075,4099,
142,213,271,334,999,1075,1736,2001,2079,2285,3159,3173,4215,4239,
44,50,67,168,724,975,1130,1242,2051,2173,2210,2742,3266,3290,
22,104,176,325,754,1079,1419,1722,1834,2395,2914,3216,3970,3994,
89,127,163,319,689,887,1588,1899,1967,2823,2989,3047,4103,4127,
27,38,91,580,595,1029,1300,1524,2109,2240,2816,3189,4245,4269,
24,69,115,145,235,718,1315,1375,2105,2395,2604,2666,3451,3475,
102,203,210,250,290,520,1290,1323,2151,2319,2370,2800,3426,3450,
54,111,242,268,712,886,1091,1127,1191,2271,2419,2586,3327,3351,
150,152,177,284,347,452,1220,1459,1532,2612,2856,2909,3668,3692,
46,118,299,312,466,852,1546,1852,2090,2307,2626,3067,3682,3706,
15,61,110,206,225,531,1611,1956,2029,2367,2691,2884,3747,3771,
21,142,266,308,440,700,1195,1780,1932,2214,2498,2860,3916,3940,
115,187,260,382,445,630,1462,1644,2081,2463,2542,3014,3598,3622,
75,137,149,329,675,873,1598,1909,1953,2809,2999,3033,4089,4113,
17,138,151,557,565,877,1326,1554,1645,2566,2617,2725,3781,3805,
121,128,135,238,730,790,1215,1771,1858,2264,2295,3159,3351,3375,
28,91,187,222,958,975,1108,1488,1979,2188,2721,3112,3244,3268,
55,188,289,827,833,906,1414,1470,1913,2535,2626,2993,4049,4073,
72,155,158,233,402,861,1482,2037,2062,2187,2562,2740,3618,3642,
24,96,301,314,468,854,1548,1854,2092,2309,2628,3069,3684,3708,
120,215,273,312,1001,1077,1738,2003,2081,2287,3161,3175,4217,4241,
14,66,75,159,250,757,1094,1435,1659,2174,2265,3044,3254,4309,
30,218,302,329,350,889,1302,1827,1969,2438,3049,3199,4105,4129,
34,65,83,210,423,791,1081,1683,1871,2875,2951,3063,4007,4031,
35,74,170,229,941,982,1115,1495,1986,2195,2728,3119,3251,3275,
31,103,308,321,475,861,1555,1861,2099,2316,2635,3052,3691,3715,
2,123,160,566,574,886,1335,1539,1654,2551,2626,2734,3790,3814,
20,185,252,472,770,951,1184,1996,2031,2426,2674,3111,4167,4191,
18,57,293,306,320,765,1267,1386,1845,2173,2466,2508,3522,3546,
31,52,98,152,218,701,1298,1382,2088,2378,2611,2673,3434,3458,
202,234,276,534,604,1021,1684,1896,1954,2210,2764,2840,3820,3844,
56,73,74,416,680,942,1496,1668,2116,2469,2576,3118,3632,3656,
43,190,306,374,1037,1067,1451,1815,2147,2253,3164,3227,4283,4307,
10,178,352,358,600,641,1396,1612,1721,2801,2889,3084,3857,3881,
131,202,284,323,988,1064,1749,2014,2068,2298,3148,3186,4204,4228,
132,206,243,489,659,930,1108,1569,1778,2649,2731,3168,3705,3729,
10,175,242,462,784,941,1198,2010,2021,2440,2664,3101,4157,4181,
181,260,351,516,795,918,1550,1998,2118,3021,3078,3125,4134,4158,
211,219,285,543,613,1030,1693,1905,1963,2219,2773,2849,3829,3853,
6,127,275,293,449,709,1180,1789,1941,2223,2507,2869,3925,3949,
28,100,305,318,472,858,1552,1858,2096,2313,2632,3049,3688,3712,
34,106,311,324,478,840,1558,1864,2102,2319,2638,3055,3694,3718,
181,236,319,336,477,802,1129,1261,1606,2341,2599,2954,3397,3421,
130,204,241,487,657,928,1106,1567,1776,2647,2729,3190,3703,3727,
34,58,101,265,405,510,1362,1590,1988,2483,2644,2670,3726,3750,
41,105,234,261,300,322,1341,1522,1885,2396,2405,2421,3477,3501,
4,67,292,303,330,751,1253,1372,1831,2183,2452,2518,3508,3532,
244,342,353,605,691,1053,1724,1771,1816,2711,2851,3092,3907,3931,
99,200,207,247,311,517,1287,1320,2148,2316,2367,2797,3423,3447,
39,103,232,259,298,320,1339,1520,1883,2394,2403,2419,3475,3499,
0,13,266,295,321,981,1466,1613,2061,2483,2918,3141,4197,4221,
130,157,193,217,299,387,1167,1237,2155,2317,2354,2544,3373,3397,
249,346,355,810,909,1008,1261,1574,1890,2286,2970,3127,4026,4050,
40,112,293,330,460,846,1540,1870,2108,2325,2620,3061,3676,3700,
34,57,64,182,738,965,1144,1232,2041,2163,2224,2756,3280,3304,
103,204,211,251,291,521,1291,1324,2152,2320,2371,2801,3427,3451,
27,49,112,279,993,1046,1748,1789,2126,2770,2778,3206,4262,4286,
62,171,296,816,834,889,1397,1477,1896,2542,2633,2976,4032,4056,
63,172,297,817,835,890,1398,1478,1897,2543,2634,2977,4033,4057,
186,217,324,341,458,807,1134,1266,1587,2346,2604,2959,3402,3426,
47,71,114,278,394,523,1351,1603,1977,2472,2657,2683,3739,3763,
258,343,356,619,681,1043,1714,1761,1806,2701,2841,3082,3897,3921,
141,215,252,498,668,915,1117,1578,1787,2658,2716,3177,3714,3738,
94,149,164,251,497,728,1567,1685,1808,2197,2888,3033,3944,3968,
99,244,287,323,329,992,1273,1409,1634,2489,2578,2641,3545,3569,
31,42,95,584,599,1009,1304,1528,2089,2244,2820,3169,4225,4249,
13,134,282,300,432,716,1187,1796,1924,2230,2514,2876,3932,3956,
155,157,182,265,352,433,1201,1440,1513,2593,2861,2914,3649,3673,
45,51,68,169,725,976,1131,1243,2052,2174,2211,2743,3267,3291,
22,190,340,346,612,629,1408,1624,1709,2789,2901,3072,3845,3869,
4,226,285,589,650,927,1669,1883,1924,2749,2986,3198,3805,3829,
21,67,116,212,231,537,1617,1962,2035,2373,2697,2890,3753,3777,
74,97,294,330,336,541,1227,1416,1505,2496,2529,2786,3552,3576,
142,145,205,229,311,399,1155,1225,2143,2305,2366,2556,3361,3385,
45,168,308,376,1039,1069,1453,1817,2149,2255,3166,3229,4285,4309,
32,54,117,284,998,1051,1729,1794,2131,2775,2783,3211,4267,4291,
81,143,155,335,681,879,1604,1915,1959,2815,2981,3039,4095,4119,
252,337,350,613,675,1037,1708,1755,1800,2695,2835,3076,3891,3915,
246,343,352,807,906,1029,1258,1571,1887,2283,2967,3124,4023,4047,
13,178,245,465,787,944,1177,2013,2024,2443,2667,3104,4160,4184,
152,206,220,496,665,829,1131,1745,1768,2338,2825,2843,3881,3905,
90,128,164,320,690,864,1589,1900,1944,2824,2990,3024,4080,4104,
44,51,93,196,409,777,1091,1693,1857,2861,2937,3049,3993,4017,
8,19,285,290,316,976,1485,1608,2056,2478,2913,3136,4192,4216,
1,122,270,288,444,704,1199,1784,1936,2218,2502,2864,3920,3944,
13,65,74,158,249,756,1093,1434,1658,2173,2264,3043,3253,4308,
5,51,100,196,239,545,1625,1946,2019,2357,2705,2898,3761,3785,
46,85,181,216,952,969,1126,1506,1973,2206,2715,3106,3262,3286,
1,14,267,296,322,982,1467,1614,2062,2484,2919,3142,4198,4222,
201,233,275,533,603,1020,1683,1919,1953,2209,2763,2839,3819,3843,
253,338,351,614,676,1038,1709,1756,1801,2696,2836,3077,3892,3916,
133,207,244,490,660,931,1109,1570,1779,2650,2732,3169,3706,3730,
1,190,257,477,775,956,1189,2001,2036,2431,2679,3116,4172,4196,
32,45,85,589,598,1023,1318,1518,2103,2234,2810,3183,4239,4263,
91,129,165,321,691,865,1590,1901,1945,2825,2991,3025,4081,4105,
46,68,107,274,988,1041,1743,1784,2121,2765,2773,3201,4257,4281,
41,113,294,331,461,847,1541,1871,2109,2326,2621,3062,3677,3701,
25,49,116,280,396,525,1353,1605,1979,2474,2659,2685,3741,3765,
57,190,291,829,835,908,1392,1472,1915,2537,2628,2995,4051,4075,
37,184,300,368,1055,1061,1445,1809,2141,2247,3158,3221,4277,4301,
56,189,290,828,834,907,1415,1471,1914,2536,2627,2994,4050,4074,
19,71,80,164,255,762,1099,1416,1664,2179,2270,3025,3259,4314,
0,121,158,564,572,884,1333,1537,1652,2549,2624,2732,3788,3812,
10,56,105,201,220,550,1630,1951,2024,2362,2710,2903,3766,3790,
146,148,173,280,343,448,1216,1455,1528,2608,2876,2905,3664,3688,
96,197,204,244,308,514,1284,1341,2145,2313,2364,2794,3420,3444,
75,145,154,256,502,733,1572,1690,1813,2202,2893,3038,3949,3973,
47,68,114,144,234,717,1314,1374,2104,2394,2603,2665,3450,3474,
72,119,292,328,358,539,1225,1438,1503,2518,2527,2784,3574,3598,
6,58,91,151,242,749,1086,1427,1675,2166,2257,3036,3246,4301,
183,262,353,518,797,920,1552,2000,2120,3023,3080,3127,4136,4160,
24,54,71,172,728,979,1134,1246,2055,2177,2214,2746,3270,3294,
173,228,335,352,469,794,1145,1253,1598,2333,2615,2970,3389,3413,
47,170,310,378,1041,1071,1455,1819,2151,2233,3144,3231,4287,4311,
13,235,270,598,659,912,1678,1892,1933,2758,2995,3207,3814,3838,
73,152,167,254,500,731,1570,1688,1811,2200,2891,3036,3947,3971,
19,184,251,471,769,950,1183,1995,2030,2425,2673,3110,4166,4190,
69,86,87,429,693,955,1509,1657,2129,2458,2589,3107,3645,3669,
42,81,177,236,948,965,1122,1502,1969,2202,2735,3102,3258,3282,
45,117,298,335,465,851,1545,1851,2089,2306,2625,3066,3681,3705,
72,134,146,326,672,870,1595,1906,1950,2830,2996,3030,4086,4110,
46,70,113,277,393,522,1350,1602,1976,2495,2656,2682,3738,3762,
125,152,212,236,294,406,1162,1232,2150,2312,2373,2563,3368,3392,
20,141,154,560,568,880,1329,1557,1648,2545,2620,2728,3784,3808,
41,65,108,272,388,517,1345,1597,1971,2490,2651,2677,3733,3757,
131,205,242,488,658,929,1107,1568,1777,2648,2730,3191,3704,3728,
156,158,183,266,353,434,1202,1441,1514,2594,2862,2915,3650,3674,
118,263,282,318,324,987,1292,1404,1653,2484,2573,2660,3540,3564,
84,154,163,241,487,742,1581,1699,1822,2187,2902,3047,3958,3982,
7,128,276,294,450,710,1181,1790,1942,2224,2508,2870,3926,3950,
14,53,289,302,316,761,1263,1382,1841,2169,2462,2504,3518,3542,
122,129,139,232,724,784,1209,1765,1852,2258,2289,3153,3345,3369,
124,151,211,235,293,405,1161,1231,2149,2311,2372,2562,3367,3391,
193,225,267,549,619,1012,1699,1911,1945,2225,2779,2855,3835,3859,
120,194,255,501,671,918,1120,1581,1790,2661,2719,3180,3717,3741,
11,125,213,269,363,557,1349,1359,1385,2348,2429,2949,3485,3509,
94,153,156,231,400,859,1480,2035,2060,2185,2560,2738,3616,3640,
25,172,288,380,1043,1073,1457,1821,2153,2235,3146,3233,4289,4313,
178,257,348,513,792,915,1547,1995,2115,3018,3075,3122,4131,4155,
14,60,109,205,224,530,1610,1955,2028,2366,2690,2883,3746,3770,
259,344,357,620,682,1044,1715,1762,1807,2702,2842,3083,3898,3922,
13,134,147,553,561,873,1322,1550,1641,2562,2637,2721,3777,3801,
263,336,345,800,899,1022,1251,1564,1880,2300,2960,3141,4016,4040,
43,82,178,237,949,966,1123,1503,1970,2203,2712,3103,3259,3283,
107,252,271,313,331,1000,1281,1393,1642,2473,2586,2649,3529,3553,
29,53,96,284,400,505,1357,1585,1983,2478,2663,2665,3721,3745,
23,62,298,311,325,746,1248,1391,1826,2178,2471,2513,3527,3551,
151,153,178,285,348,453,1221,1460,1533,2613,2857,2910,3669,3693,
102,247,266,326,332,995,1276,1412,1637,2492,2581,2644,3548,3572,
3,14,280,309,335,971,1480,1627,2051,2473,2908,3131,4187,4211,
165,195,233,485,654,818,1144,1734,1757,2351,2814,2832,3870,3894,
5,111,183,332,761,1062,1426,1705,1841,2378,2921,3223,3977,4001,
118,190,263,361,448,633,1441,1647,2084,2466,2521,3017,3577,3601,
81,151,160,262,484,739,1578,1696,1819,2184,2899,3044,3955,3979,
2,15,268,297,323,983,1468,1615,2063,2485,2920,3143,4199,4223,
130,201,283,322,987,1063,1748,2013,2067,2297,3147,3185,4203,4227,
113,258,277,313,319,1006,1287,1399,1648,2479,2568,2655,3535,3559,
41,80,176,235,947,964,1121,1501,1968,2201,2734,3101,3257,3281,
97,198,205,245,309,515,1285,1342,2146,2314,2365,2795,3421,3445,
24,37,77,581,590,1015,1310,1534,2095,2250,2826,3175,4231,4255,
126,133,140,219,735,771,1220,1752,1863,2269,2300,3164,3356,3380,
213,221,287,545,615,1008,1695,1907,1965,2221,2775,2851,3831,3855,
102,174,247,369,432,641,1449,1655,2068,2450,2529,3001,3585,3609,
108,192,209,256,296,526,1272,1329,2157,2325,2352,2806,3408,3432,
125,199,260,482,652,923,1125,1562,1795,2642,2724,3185,3698,3722,
129,203,240,486,656,927,1105,1566,1799,2646,2728,3189,3702,3726,
5,143,207,287,381,575,1353,1367,1379,2342,2447,2943,3503,3527,
46,52,69,170,726,977,1132,1244,2053,2175,2212,2744,3268,3292,
29,51,114,281,995,1048,1750,1791,2128,2772,2780,3208,4264,4288,
12,23,265,294,320,980,1465,1612,2060,2482,2917,3140,4196,4220,
151,205,219,495,664,828,1130,1744,1767,2337,2824,2842,3880,3904,
41,48,90,193,430,774,1088,1690,1854,2858,2934,3070,3990,4014,
78,148,157,259,481,736,1575,1693,1816,2205,2896,3041,3952,3976,
196,228,270,528,622,1015,1702,1914,1948,2228,2782,2834,3838,3862,
177,232,315,356,473,798,1149,1257,1602,2337,2595,2974,3393,3417,
73,156,159,234,403,862,1483,2038,2063,2188,2563,2741,3619,3643,
39,111,292,329,459,845,1539,1869,2107,2324,2619,3060,3675,3699,
27,90,186,221,957,974,1107,1511,1978,2187,2720,3111,3243,3267,
64,97,252,278,698,872,1101,1113,1177,2257,2405,2572,3313,3337,
174,253,344,509,812,935,1543,2015,2135,3014,3095,3142,4151,4175,
24,55,73,200,413,781,1095,1697,1861,2865,2941,3053,3997,4021,
2,65,290,301,328,749,1251,1370,1829,2181,2450,2516,3506,3530,
52,185,310,824,830,903,1411,1467,1910,2532,2623,2990,4046,4070,
53,94,95,413,677,939,1493,1665,2113,2466,2573,3115,3629,3653,
25,113,218,245,308,330,1325,1530,1893,2380,2405,2413,3461,3485,
178,233,316,357,474,799,1150,1258,1603,2338,2596,2975,3394,3418,
11,50,299,310,313,758,1260,1379,1838,2166,2459,2501,3515,3539,
72,141,268,347,641,848,1281,1928,2067,2701,2938,3008,4064,4088,
34,181,297,365,1052,1058,1442,1806,2138,2244,3155,3218,4274,4298,
103,175,248,370,433,642,1450,1632,2069,2451,2530,3002,3586,3610,
1,64,289,300,327,748,1250,1369,1828,2180,2449,2515,3505,3529,
261,346,359,622,684,1046,1717,1764,1809,2704,2844,3085,3900,3924,
89,112,309,321,351,532,1242,1431,1496,2511,2520,2801,3567,3591,
76,138,150,330,676,874,1599,1910,1954,2810,2976,3034,4090,4114,
80,125,276,355,625,856,1289,1936,2075,2709,2946,3016,4072,4096,
28,216,300,327,348,911,1300,1825,1991,2436,3071,3197,4127,4151,
10,232,267,595,656,933,1675,1889,1930,2755,2992,3204,3811,3835,
189,244,359,524,803,926,1558,2006,2126,3005,3086,3133,4142,4166,
47,86,182,217,953,970,1127,1507,1974,2207,2716,3107,3263,3287,
121,192,274,313,1002,1078,1739,2004,2082,2288,3162,3176,4218,4242,
42,114,295,332,462,848,1542,1848,2110,2327,2622,3063,3678,3702,
133,160,196,220,302,390,1170,1240,2158,2320,2357,2547,3376,3400,
3,225,284,588,649,926,1668,1882,1923,2748,2985,3197,3804,3828,
116,261,280,316,322,985,1290,1402,1651,2482,2571,2658,3538,3562,
71,88,89,431,695,957,1511,1659,2131,2460,2591,3109,3647,3671,
159,161,186,269,356,437,1205,1444,1517,2597,2865,2918,3653,3677,
79,102,299,335,341,546,1232,1421,1510,2501,2534,2791,3557,3581,
127,154,214,238,296,384,1164,1234,2152,2314,2375,2565,3370,3394,
87,125,161,317,687,885,1586,1897,1965,2821,2987,3045,4101,4125,
38,110,291,328,458,844,1538,1868,2106,2323,2618,3059,3674,3698,
29,40,93,582,597,1031,1302,1526,2111,2242,2818,3191,4247,4271,
46,67,113,167,233,716,1313,1373,2103,2393,2602,2664,3449,3473,
2,224,283,587,648,925,1667,1881,1922,2747,2984,3196,3803,3827,
136,207,265,328,993,1069,1730,1995,2073,2303,3153,3191,4209,4233,
91,114,311,323,353,534,1244,1433,1498,2513,2522,2803,3569,3593,
82,134,186,205,214,415,1162,1164,1223,2242,2965,3234,3298,3322,
2,191,258,478,776,957,1190,2002,2037,2432,2680,3117,4173,4197,
0,63,288,299,326,747,1249,1368,1827,2179,2448,2514,3504,3528,
206,238,280,538,608,1025,1688,1900,1958,2214,2768,2844,3824,3848,
248,346,357,609,695,1033,1704,1775,1820,2691,2855,3072,3911,3935,
33,46,86,590,599,1024,1319,1519,2104,2235,2811,3184,4240,4264,
0,106,178,327,756,1057,1421,1724,1836,2397,2916,3218,3972,3996,
157,211,225,501,670,834,1136,1750,1773,2343,2830,2848,3886,3910,
29,117,222,249,288,334,1329,1534,1873,2384,2409,2417,3465,3489,
36,59,66,184,740,967,1146,1234,2043,2165,2226,2758,3282,3306,
91,136,287,342,636,843,1276,1923,2086,2696,2933,3003,4059,4083,
163,165,190,273,336,441,1209,1448,1521,2601,2869,2922,3657,3681,
139,210,268,331,996,1072,1733,1998,2076,2282,3156,3170,4212,4236,
31,119,224,251,290,312,1331,1512,1875,2386,2411,2419,3467,3491,
197,229,271,529,623,1016,1703,1915,1949,2229,2783,2835,3839,3863,
195,227,269,551,621,1014,1701,1913,1947,2227,2781,2833,3837,3861,
121,128,138,231,723,783,1208,1764,1851,2257,2288,3152,3344,3368,
125,132,139,218,734,770,1219,1775,1862,2268,2299,3163,3355,3379,
77,147,156,258,480,735,1574,1692,1815,2204,2895,3040,3951,3975,
9,123,211,267,361,555,1347,1357,1383,2346,2427,2947,3483,3507,
33,105,310,323,477,863,1557,1863,2101,2318,2637,3054,3693,3717,
90,145,160,247,493,724,1563,1681,1804,2193,2884,3029,3940,3964,
179,234,317,358,475,800,1151,1259,1604,2339,2597,2952,3395,3419,
55,72,73,415,679,941,1495,1667,2115,2468,2575,3117,3631,3655,
4,172,346,352,618,635,1414,1630,1715,2795,2883,3078,3851,3875,
179,258,349,514,793,916,1548,1996,2116,3019,3076,3123,4132,4156,
8,230,265,593,654,931,1673,1887,1928,2753,2990,3202,3809,3833,
11,117,189,314,767,1068,1432,1711,1847,2384,2927,3229,3983,4007,
45,66,112,166,232,715,1312,1372,2102,2392,2601,2687,3448,3472,
43,107,236,263,302,324,1343,1524,1887,2398,2407,2423,3479,3503,
160,162,187,270,357,438,1206,1445,1518,2598,2866,2919,3654,3678,
31,55,98,286,402,507,1359,1587,1985,2480,2641,2667,3723,3747,
32,56,99,287,403,508,1360,1588,1986,2481,2642,2668,3724,3748,
68,177,302,816,822,895,1403,1483,1902,2524,2639,2982,4038,4062,
84,146,167,221,390,849,1470,2025,2050,2199,2550,2752,3606,3630,
4,125,273,291,447,707,1178,1787,1939,2221,2505,2867,3923,3947,
153,155,180,287,350,455,1223,1462,1535,2615,2859,2912,3671,3695,
133,204,286,325,990,1066,1751,1992,2070,2300,3150,3188,4206,4230,
145,199,237,489,658,822,1148,1738,1761,2331,2818,2836,3874,3898,
126,200,261,483,653,924,1126,1563,1796,2643,2725,3186,3699,3723,
20,102,174,323,752,1077,1417,1720,1832,2393,2912,3238,3968,3992,
40,64,107,271,387,516,1344,1596,1970,2489,2650,2676,3732,3756,
5,126,163,553,569,865,1338,1542,1633,2554,2629,2713,3769,3793,
80,132,184,203,212,413,1160,1162,1221,2240,2963,3232,3296,3320,
23,120,157,563,571,883,1332,1536,1651,2548,2623,2731,3787,3811,
10,131,144,558,574,870,1343,1547,1638,2559,2634,2718,3774,3798,
46,53,95,198,411,779,1093,1695,1859,2863,2939,3051,3995,4019,
158,160,185,268,355,436,1204,1443,1516,2596,2864,2917,3652,3676,
118,195,202,242,306,512,1282,1339,2143,2311,2362,2792,3418,3442,
8,60,93,153,244,751,1088,1429,1677,2168,2259,3038,3248,4303,
32,179,295,363,1050,1056,1440,1804,2136,2242,3153,3216,4272,4296,
7,175,349,355,621,638,1393,1609,1718,2798,2886,3081,3854,3878,
4,17,270,299,325,961,1470,1617,2041,2487,2922,3121,4177,4201,
129,200,282,321,986,1062,1747,2012,2066,2296,3146,3184,4202,4226,
95,123,175,194,203,428,1153,1175,1212,2255,2954,3223,3311,3335,
29,101,306,319,473,859,1553,1859,2097,2314,2633,3050,3689,3713,
129,156,192,216,298,386,1166,1236,2154,2316,2353,2567,3372,3396,
115,260,279,315,321,984,1289,1401,1650,2481,2570,2657,3537,3561,
27,40,80,584,593,1018,1313,1513,2098,2253,2829,3178,4234,4258,
43,67,110,274,390,519,1347,1599,1973,2492,2653,2679,3735,3759,
22,61,297,310,324,745,1271,1390,1825,2177,2470,2512,3526,3550,
49,106,261,287,707,881,1086,1122,1186,2266,2414,2581,3322,3346,
191,246,337,526,805,928,1536,2008,2128,3007,3088,3135,4144,4168,
11,179,353,359,601,642,1397,1613,1722,2802,2890,3085,3858,3882,
77,160,163,238,407,842,1487,2018,2043,2192,2567,2745,3623,3647,
21,60,296,309,323,744,1270,1389,1824,2176,2469,2511,3525,3549,
93,152,155,230,399,858,1479,2034,2059,2184,2559,2737,3615,3639,
40,104,233,260,299,321,1340,1521,1884,2395,2404,2420,3476,3500,
3,55,88,148,263,746,1083,1424,1672,2163,2278,3033,3243,4298,
26,71,117,147,237,696,1317,1377,2107,2397,2606,2668,3453,3477,
0,121,269,311,443,703,1198,1783,1935,2217,2501,2863,3919,3943,
128,155,215,239,297,385,1165,1235,2153,2315,2352,2566,3371,3395,
27,48,118,148,238,697,1318,1378,2108,2398,2607,2669,3454,3478,
96,241,284,320,326,989,1294,1406,1655,2486,2575,2662,3542,3566,
87,139,191,195,210,420,1167,1169,1204,2247,2970,3239,3303,3327,
240,337,346,801,900,1023,1252,1565,1881,2301,2961,3142,4017,4041,
80,150,159,261,483,738,1577,1695,1818,2207,2898,3043,3954,3978,
256,338,353,793,892,1015,1268,1581,1873,2293,2953,3134,4009,4033,
19,133,197,277,371,565,1357,1367,1369,2332,2437,2933,3493,3517,
9,231,266,594,655,932,1674,1888,1929,2754,2991,3203,3810,3834,
104,249,268,328,334,997,1278,1414,1639,2494,2583,2646,3550,3574,
40,71,89,192,429,773,1087,1689,1853,2857,2933,3069,3989,4013,
180,259,350,515,794,917,1549,1997,2117,3020,3077,3124,4133,4157,
137,208,266,329,994,1070,1731,1996,2074,2280,3154,3168,4210,4234,
18,183,250,470,768,949,1182,1994,2029,2424,2672,3109,4165,4189,
93,131,167,323,693,867,1592,1903,1947,2827,2993,3027,4083,4107,
41,62,108,162,228,711,1308,1368,2098,2388,2597,2683,3444,3468,
4,56,89,149,240,747,1084,1425,1673,2164,2279,3034,3244,4299,
80,103,300,312,342,547,1233,1422,1511,2502,2535,2792,3558,3582,
95,154,157,232,401,860,1481,2036,2061,2186,2561,2739,3617,3641,
73,125,177,196,205,430,1153,1155,1214,2233,2956,3225,3289,3313,
139,166,202,226,308,396,1152,1246,2140,2326,2363,2553,3382,3406,
21,135,199,279,373,567,1345,1359,1371,2334,2439,2935,3495,3519,
46,110,239,242,305,327,1322,1527,1890,2377,2402,2410,3458,3482,
10,62,95,155,246,753,1090,1431,1679,2170,2261,3040,3250,4305,
164,194,232,484,653,817,1143,1733,1756,2350,2813,2855,3869,3893,
88,158,167,245,491,722,1561,1703,1802,2191,2882,3027,3938,3962,
35,56,102,156,222,705,1302,1386,2092,2382,2615,2677,3438,3462,
95,133,145,325,695,869,1594,1905,1949,2829,2995,3029,4085,4109,
112,196,213,260,300,506,1276,1333,2137,2305,2356,2786,3412,3436,
21,103,175,324,753,1078,1418,1721,1833,2394,2913,3239,3969,3993,
16,137,150,556,564,876,1325,1553,1644,2565,2616,2724,3780,3804,
147,149,174,281,344,449,1217,1456,1529,2609,2877,2906,3665,3689,
29,217,301,328,349,888,1301,1826,1968,2437,3048,3198,4104,4128,
23,51,84,144,259,766,1103,1420,1668,2183,2274,3029,3263,4318,
122,149,209,233,291,403,1159,1229,2147,2309,2370,2560,3365,3389,
89,141,169,197,212,422,1169,1171,1206,2249,2972,3217,3305,3329,
263,337,348,600,686,1048,1719,1766,1811,2706,2846,3087,3902,3926,
1,223,282,586,671,924,1666,1880,1921,2746,2983,3195,3802,3826,
12,180,336,354,602,643,1398,1614,1723,2803,2891,3086,3859,3883,
18,70,79,163,254,761,1098,1439,1663,2178,2269,3024,3258,4313,
101,246,265,325,331,994,1275,1411,1636,2491,2580,2643,3547,3571,
24,171,311,379,1042,1072,1456,1820,2152,2234,3145,3232,4288,4312,
50,183,308,822,828,901,1409,1465,1908,2530,2621,2988,4044,4068,
13,181,337,355,603,644,1399,1615,1724,2804,2892,3087,3860,3884,
84,107,304,316,346,551,1237,1426,1491,2506,2539,2796,3562,3586,
94,132,144,324,694,868,1593,1904,1948,2828,2994,3028,4084,4108,
24,112,217,244,307,329,1324,1529,1892,2379,2404,2412,3460,3484,
19,187,337,343,609,626,1405,1621,1706,2786,2898,3093,3842,3866,
148,150,175,282,345,450,1218,1457,1530,2610,2878,2907,3666,3690,
205,237,279,537,607,1024,1687,1899,1957,2213,2767,2843,3823,3847,
165,167,168,275,338,443,1211,1450,1523,2603,2871,2924,3659,3683,
90,135,286,341,635,842,1275,1922,2085,2695,2932,3002,4058,4082,
7,18,284,289,315,975,1484,1631,2055,2477,2912,3135,4191,4215,
45,67,106,273,987,1040,1742,1783,2120,2764,2772,3200,4256,4280,
173,252,343,508,811,934,1542,2014,2134,3013,3094,3141,4150,4174,
113,197,214,261,301,507,1277,1334,2138,2306,2357,2787,3413,3437,
74,157,160,235,404,863,1484,2039,2040,2189,2564,2742,3620,3644,
121,131,138,224,740,776,1201,1757,1868,2274,2281,3145,3337,3361,
67,176,301,821,839,894,1402,1482,1901,2523,2638,2981,4037,4061,
91,146,161,248,494,725,1564,1682,1805,2194,2885,3030,3941,3965,
90,149,152,227,396,855,1476,2031,2056,2205,2556,2758,3612,3636,
37,101,230,257,296,318,1337,1518,1881,2392,2401,2417,3473,3497,
10,124,212,268,362,556,1348,1358,1384,2347,2428,2948,3484,3508,
25,56,74,201,414,782,1096,1698,1862,2866,2942,3054,3998,4022,
15,67,76,160,251,758,1095,1436,1660,2175,2266,3045,3255,4310,
17,185,341,359,607,624,1403,1619,1704,2784,2896,3091,3840,3864,
41,63,102,269,1007,1036,1738,1779,2116,2760,2768,3196,4252,4276,
2,170,344,350,616,633,1412,1628,1713,2793,2881,3076,3849,3873,
47,53,70,171,727,978,1133,1245,2054,2176,2213,2745,3269,3293,
7,20,273,302,328,964,1473,1620,2044,2490,2925,3124,4180,4204,
87,157,166,244,490,721,1560,1702,1801,2190,2881,3026,3937,3961,
73,142,269,348,642,849,1282,1929,2068,2702,2939,3009,4065,4089,
251,336,349,612,674,1036,1707,1754,1823,2694,2834,3075,3890,3914,
53,186,311,825,831,904,1412,1468,1911,2533,2624,2991,4047,4071,
84,129,280,359,629,860,1293,1940,2079,2689,2950,3020,4076,4100,
207,239,281,539,609,1026,1689,1901,1959,2215,2769,2845,3825,3849,
115,192,199,263,303,509,1279,1336,2140,2308,2359,2789,3415,3439,
26,37,90,579,594,1028,1299,1523,2108,2239,2815,3188,4244,4268,
7,113,185,334,763,1064,1428,1707,1843,2380,2923,3225,3979,4003,
64,173,298,818,836,891,1399,1479,1898,2520,2635,2978,4034,4058,
48,181,306,820,826,899,1407,1487,1906,2528,2619,2986,4042,4066,
99,171,244,366,453,638,1446,1652,2065,2471,2526,3022,3582,3606,
5,68,293,304,331,752,1254,1373,1832,2160,2453,2519,3509,3533,
66,83,84,426,690,952,1506,1678,2126,2455,2586,3104,3642,3666,
103,248,267,327,333,996,1277,1413,1638,2493,2582,2645,3549,3573,
11,233,268,596,657,934,1676,1890,1931,2756,2993,3205,3812,3836,
106,251,270,312,330,999,1280,1392,1641,2472,2585,2648,3528,3552,
70,179,304,818,824,897,1405,1485,1904,2526,2617,2984,4040,4064,
8,54,103,199,218,548,1628,1949,2022,2360,2708,2901,3764,3788,
44,68,111,275,391,520,1348,1600,1974,2493,2654,2680,3736,3760,
33,221,305,332,353,892,1305,1830,1972,2441,3052,3202,4108,4132,
61,78,79,421,685,947,1501,1673,2121,2450,2581,3099,3637,3661,
15,136,284,302,434,718,1189,1798,1926,2208,2516,2878,3934,3958,
126,197,279,318,1007,1059,1744,2009,2087,2293,3167,3181,4223,4247,
42,230,290,317,338,901,1314,1839,1981,2426,3061,3211,4117,4141,
78,130,182,201,210,411,1158,1160,1219,2238,2961,3230,3294,3318,
16,98,170,319,748,1073,1437,1716,1828,2389,2908,3234,3964,3988,
143,146,206,230,288,400,1156,1226,2144,2306,2367,2557,3362,3386,
185,216,323,340,457,806,1133,1265,1586,2345,2603,2958,3401,3425,
43,49,66,191,723,974,1129,1241,2050,2172,2209,2741,3265,3289,
36,108,289,326,456,842,1536,1866,2104,2321,2616,3057,3672,3696,
0,222,281,585,670,923,1665,1879,1920,2745,2982,3194,3801,3825,
176,231,314,355,472,797,1148,1256,1601,2336,2594,2973,3392,3416,
39,60,106,160,226,709,1306,1390,2096,2386,2595,2681,3442,3466,
26,57,75,202,415,783,1097,1699,1863,2867,2943,3055,3999,4023,
15,97,169,318,747,1072,1436,1715,1827,2388,2907,3233,3963,3987,
16,130,194,274,368,562,1354,1364,1390,2329,2434,2930,3490,3514,
1,71,96,192,235,541,1621,1966,2039,2353,2701,2894,3757,3781,
22,136,200,280,374,568,1346,1360,1372,2335,2440,2936,3496,3520,
257,342,355,618,680,1042,1713,1760,1805,2700,2840,3081,3896,3920,
44,66,105,272,986,1039,1741,1782,2119,2763,2771,3199,4255,4279,
33,55,118,285,999,1052,1730,1795,2132,2760,2776,3212,4268,4292,
7,229,264,592,653,930,1672,1886,1927,2752,2989,3201,3808,3832,
19,58,294,307,321,766,1268,1387,1846,2174,2467,2509,3523,3547,
65,174,299,819,837,892,1400,1480,1899,2521,2636,2979,4035,4059,
35,107,288,325,479,841,1559,1865,2103,2320,2639,3056,3695,3719,
10,21,287,292,318,978,1487,1610,2058,2480,2915,3138,4194,4218,
22,68,117,213,232,538,1618,1963,2036,2374,2698,2891,3754,3778,
174,229,312,353,470,795,1146,1254,1599,2334,2592,2971,3390,3414,
140,167,203,227,309,397,1153,1247,2141,2327,2364,2554,3383,3407,
21,219,278,582,667,920,1662,1876,1941,2742,2979,3215,3798,3822,
35,182,298,366,1053,1059,1443,1807,2139,2245,3156,3219,4275,4299,
126,136,143,229,721,781,1206,1762,1849,2279,2286,3150,3342,3366,
21,49,82,166,257,764,1101,1418,1666,2181,2272,3027,3261,4316,
2,48,97,193,236,542,1622,1967,2016,2354,2702,2895,3758,3782,
119,196,203,243,307,513,1283,1340,2144,2312,2363,2793,3419,3443,
8,122,210,266,360,554,1346,1356,1382,2345,2426,2946,3482,3506,
42,189,305,373,1036,1066,1450,1814,2146,2252,3163,3226,4282,4306,
34,47,87,576,591,1025,1296,1520,2105,2236,2812,3185,4241,4265,
92,115,288,324,354,535,1245,1434,1499,2514,2523,2804,3570,3594,
13,127,215,271,365,559,1351,1361,1387,2350,2431,2951,3487,3511,
53,110,241,267,711,885,1090,1126,1190,2270,2418,2585,3326,3350,
77,129,181,200,209,410,1157,1159,1218,2237,2960,3229,3293,3317,
35,58,65,183,739,966,1145,1233,2042,2164,2225,2757,3281,3305,
259,341,356,796,895,1018,1271,1560,1876,2296,2956,3137,4012,4036,
93,148,163,250,496,727,1566,1684,1807,2196,2887,3032,3943,3967,
84,122,158,314,684,882,1607,1918,1962,2818,2984,3042,4098,4122,
12,126,214,270,364,558,1350,1360,1386,2349,2430,2950,3486,3510,
34,56,119,286,1000,1053,1731,1796,2133,2761,2777,3213,4269,4293,
20,134,198,278,372,566,1344,1358,1370,2333,2438,2934,3494,3518,
243,340,349,804,903,1026,1255,1568,1884,2280,2964,3121,4020,4044,
15,136,149,555,563,875,1324,1552,1643,2564,2639,2723,3779,3803,
33,57,100,264,404,509,1361,1589,1987,2482,2643,2669,3725,3749,
250,348,359,611,673,1035,1706,1753,1822,2693,2833,3074,3889,3913,
91,143,171,199,214,424,1171,1173,1208,2251,2974,3219,3307,3331,
29,60,78,205,418,786,1100,1702,1866,2870,2946,3058,4002,4026,
6,120,208,264,382,552,1344,1354,1380,2343,2424,2944,3480,3504,
3,49,98,194,237,543,1623,1944,2017,2355,2703,2896,3759,3783,
61,170,295,833,839,888,1396,1476,1919,2541,2632,2999,4055,4079,
18,100,172,321,750,1075,1439,1718,1830,2391,2910,3236,3966,3990,
96,168,241,363,450,635,1443,1649,2086,2468,2523,3019,3579,3603,
253,350,359,814,889,1012,1265,1578,1894,2290,2974,3131,4030,4054,
16,62,111,207,226,532,1612,1957,2030,2368,2692,2885,3748,3772,
65,82,83,425,689,951,1505,1677,2125,2454,2585,3103,3641,3665,
37,76,172,231,943,960,1117,1497,1988,2197,2730,3097,3253,3277,
111,195,212,259,299,505,1275,1332,2136,2304,2355,2785,3411,3435,
69,102,257,283,703,877,1082,1118,1182,2262,2410,2577,3318,3342,
12,234,269,597,658,935,1677,1891,1932,2757,2994,3206,3813,3837,
17,182,249,469,791,948,1181,1993,2028,2447,2671,3108,4164,4188,
39,186,302,370,1033,1063,1447,1811,2143,2249,3160,3223,4279,4303,
18,216,275,579,664,917,1659,1873,1938,2739,2976,3212,3795,3819,
36,224,308,335,356,895,1308,1833,1975,2444,3055,3205,4111,4135,
15,180,247,467,789,946,1179,2015,2026,2445,2669,3106,4162,4186,
121,195,256,502,648,919,1121,1582,1791,2662,2720,3181,3718,3742,
161,215,229,481,650,838,1140,1730,1753,2347,2810,2852,3866,3890,
138,212,249,495,665,912,1114,1575,1784,2655,2713,3174,3711,3735,
27,115,220,247,310,332,1327,1532,1895,2382,2407,2415,3463,3487,
110,182,255,377,440,625,1457,1639,2076,2458,2537,3009,3593,3617,
38,59,105,159,225,708,1305,1389,2095,2385,2594,2680,3441,3465,
1,53,86,146,261,744,1081,1422,1670,2161,2276,3031,3241,4296,
14,96,168,317,746,1071,1435,1714,1826,2387,2906,3232,3962,3986,
20,66,115,211,230,536,1616,1961,2034,2372,2696,2889,3752,3776,
35,59,102,266,406,511,1363,1591,1989,2484,2645,2671,3727,3751,
140,214,251,497,667,914,1116,1577,1786,2657,2715,3176,3713,3737,
248,345,354,809,908,1031,1260,1573,1889,2285,2969,3126,4025,4049,
114,198,215,262,302,508,1278,1335,2139,2307,2358,2788,3414,3438,
168,223,330,347,464,813,1140,1248,1593,2328,2610,2965,3384,3408,
95,140,267,346,640,847,1280,1927,2066,2700,2937,3007,4063,4087,
117,262,281,317,323,986,1291,1403,1652,2483,2572,2659,3539,3563,
41,188,304,372,1035,1065,1449,1813,2145,2251,3162,3225,4281,4305,
63,80,81,423,687,949,1503,1675,2123,2452,2583,3101,3639,3663,
97,169,242,364,451,636,1444,1650,2087,2469,2524,3020,3580,3604,
28,52,119,283,399,504,1356,1584,1982,2477,2662,2664,3720,3744,
30,61,79,206,419,787,1101,1703,1867,2871,2947,3059,4003,4027,
112,257,276,312,318,1005,1286,1398,1647,2478,2591,2654,3534,3558,
27,58,76,203,416,784,1098,1700,1864,2868,2944,3056,4000,4024,
69,178,303,817,823,896,1404,1484,1903,2525,2616,2983,4039,4063,
245,343,354,606,692,1054,1725,1772,1817,2688,2852,3093,3908,3932,
109,193,210,257,297,527,1273,1330,2158,2326,2353,2807,3409,3433,
36,75,171,230,942,983,1116,1496,1987,2196,2729,3096,3252,3276,
68,85,86,428,692,954,1508,1656,2128,2457,2588,3106,3644,3668,
1,169,343,349,615,632,1411,1627,1712,2792,2880,3075,3848,3872,
19,140,153,559,567,879,1328,1556,1647,2544,2619,2727,3783,3807,
26,89,185,220,956,973,1106,1510,1977,2186,2719,3110,3242,3266,
44,83,179,238,950,967,1124,1504,1971,2204,2713,3104,3260,3284,
58,191,292,830,836,909,1393,1473,1916,2538,2629,2996,4052,4076,
1,139,203,283,377,571,1349,1363,1375,2338,2443,2939,3499,3523,
36,67,85,212,425,769,1083,1685,1849,2877,2929,3065,3985,4009,
112,184,257,379,442,627,1459,1641,2078,2460,2539,3011,3595,3619,
28,50,113,280,994,1047,1749,1790,2127,2771,2779,3207,4263,4287,
9,115,187,312,765,1066,1430,1709,1845,2382,2925,3227,3981,4005,
37,61,104,268,384,513,1365,1593,1991,2486,2647,2673,3729,3753,
84,136,188,192,207,417,1164,1166,1201,2244,2967,3236,3300,3324,
43,64,110,164,230,713,1310,1370,2100,2390,2599,2685,3446,3470,
124,134,141,227,743,779,1204,1760,1871,2277,2284,3148,3340,3364,
49,90,91,409,673,959,1489,1661,2133,2462,2569,3111,3625,3649,
9,61,94,154,245,752,1089,1430,1678,2169,2260,3039,3249,4304,
42,106,235,262,301,323,1342,1523,1886,2397,2406,2422,3478,3502,
176,255,346,511,814,913,1545,1993,2113,3016,3073,3120,4129,4153,
187,218,325,342,459,808,1135,1267,1588,2347,2605,2960,3403,3427,
45,233,293,320,341,904,1317,1842,1984,2429,3064,3214,4120,4144,
59,116,247,273,717,867,1096,1108,1196,2276,2400,2591,3332,3356,
15,183,339,357,605,646,1401,1617,1726,2806,2894,3089,3862,3886,
188,243,358,523,802,925,1557,2005,2125,3004,3085,3132,4141,4165,
67,100,255,281,701,875,1080,1116,1180,2260,2408,2575,3316,3340,
17,131,195,275,369,563,1355,1365,1391,2330,2435,2931,3491,3515,
26,49,56,174,730,981,1136,1224,2057,2179,2216,2748,3272,3296,
184,263,354,519,798,921,1553,2001,2121,3000,3081,3128,4137,4161,
16,181,248,468,790,947,1180,1992,2027,2446,2670,3107,4163,4187,
76,146,155,257,503,734,1573,1691,1814,2203,2894,3039,3950,3974,
40,187,303,371,1034,1064,1448,1812,2144,2250,3161,3224,4280,4304,
114,259,278,314,320,1007,1288,1400,1649,2480,2569,2656,3536,3560,
10,116,188,313,766,1067,1431,1710,1846,2383,2926,3228,3982,4006,
83,106,303,315,345,550,1236,1425,1490,2505,2538,2795,3561,3585,
134,208,245,491,661,932,1110,1571,1780,2651,2733,3170,3707,3731,
4,15,281,310,312,972,1481,1628,2052,2474,2909,3132,4188,4212,
20,218,277,581,666,919,1661,1875,1940,2741,2978,3214,3797,3821,
14,179,246,466,788,945,1178,2014,2025,2444,2668,3105,4161,4185,
6,174,348,354,620,637,1392,1608,1717,2797,2885,3080,3853,3877,
38,77,173,232,944,961,1118,1498,1989,2198,2731,3098,3254,3278,
32,104,309,322,476,862,1556,1862,2100,2317,2636,3053,3692,3716,
23,69,118,214,233,539,1619,1964,2037,2375,2699,2892,3755,3779,
106,178,251,373,436,645,1453,1635,2072,2454,2533,3005,3589,3613,
116,193,200,240,304,510,1280,1337,2141,2309,2360,2790,3416,3440,
43,115,296,333,463,849,1543,1849,2111,2304,2623,3064,3679,3703,
18,132,196,276,370,564,1356,1366,1368,2331,2436,2932,3492,3516,
31,53,116,283,997,1050,1728,1793,2130,2774,2782,3210,4266,4290,
23,221,280,584,669,922,1664,1878,1943,2744,2981,3193,3800,3824,
26,98,303,316,470,856,1550,1856,2094,2311,2630,3071,3686,3710,
120,130,137,223,739,775,1200,1756,1867,2273,2280,3144,3336,3360,
57,74,75,417,681,943,1497,1669,2117,2470,2577,3119,3633,3657,
88,140,168,196,211,421,1168,1170,1205,2248,2971,3216,3304,3328,
8,176,350,356,622,639,1394,1610,1719,2799,2887,3082,3855,3879,
38,102,231,258,297,319,1338,1519,1882,2393,2402,2418,3474,3498,
74,126,178,197,206,431,1154,1156,1215,2234,2957,3226,3290,3314,
122,196,257,503,649,920,1122,1583,1792,2663,2721,3182,3719,3743,
45,69,112,276,392,521,1349,1601,1975,2494,2655,2681,3737,3761,
194,226,268,550,620,1013,1700,1912,1946,2226,2780,2832,3836,3860,
37,109,290,327,457,843,1537,1867,2105,2322,2617,3058,3673,3697,
78,123,274,353,647,854,1287,1934,2073,2707,2944,3014,4070,4094,
104,176,249,371,434,643,1451,1633,2070,2452,2531,3003,3587,3611,
62,79,80,422,686,948,1502,1674,2122,2451,2582,3100,3638,3662,
40,61,107,161,227,710,1307,1391,2097,2387,2596,2682,3443,3467,
132,203,285,324,989,1065,1750,2015,2069,2299,3149,3187,4205,4229,
245,342,351,806,905,1028,1257,1570,1886,2282,2966,3123,4022,4046,
38,62,105,269,385,514,1366,1594,1968,2487,2648,2674,3730,3754,
124,198,259,481,651,922,1124,1561,1794,2641,2723,3184,3697,3721,
86,131,282,337,631,862,1295,1942,2081,2691,2928,3022,4078,4102,
77,100,297,333,339,544,1230,1419,1508,2499,2532,2789,3555,3579,
127,201,262,484,654,925,1127,1564,1797,2644,2726,3187,3700,3724,
74,144,153,255,501,732,1571,1689,1812,2201,2892,3037,3948,3972,
105,250,269,329,335,998,1279,1415,1640,2495,2584,2647,3551,3575,
1,107,179,328,757,1058,1422,1725,1837,2398,2917,3219,3973,3997,
5,170,261,457,779,936,1193,2005,2016,2435,2683,3096,4152,4176,
73,96,293,329,359,540,1226,1439,1504,2519,2528,2785,3575,3599,
44,65,111,165,231,714,1311,1371,2101,2391,2600,2686,3447,3471,
139,213,250,496,666,913,1115,1576,1785,2656,2714,3175,3712,3736,
51,92,93,411,675,937,1491,1663,2135,2464,2571,3113,3627,3651,
100,172,245,367,454,639,1447,1653,2066,2448,2527,3023,3583,3607,
24,48,115,279,395,524,1352,1604,1978,2473,2658,2684,3740,3764,
32,53,99,153,219,702,1299,1383,2089,2379,2612,2674,3435,3459,
42,49,91,194,431,775,1089,1691,1855,2859,2935,3071,3991,4015,
48,105,260,286,706,880,1085,1121,1185,2265,2413,2580,3321,3345,
35,66,84,211,424,768,1082,1684,1848,2876,2928,3064,3984,4008,
14,182,338,356,604,645,1400,1616,1725,2805,2893,3088,3861,3885,
242,340,351,603,689,1051,1722,1769,1814,2709,2849,3090,3905,3929,
51,184,309,823,829,902,1410,1466,1909,2531,2622,2989,4045,4069,
108,253,272,314,332,1001,1282,1394,1643,2474,2587,2650,3530,3554,
121,148,208,232,290,402,1158,1228,2146,2308,2369,2559,3364,3388,
2,54,87,147,262,745,1082,1423,1671,2162,2277,3032,3242,4297,
184,239,322,339,456,805,1132,1264,1585,2344,2602,2957,3400,3424,
192,224,266,548,618,1011,1698,1910,1944,2224,2778,2854,3834,3858,
3,168,259,479,777,958,1191,2003,2038,2433,2681,3118,4174,4198,
2,123,271,289,445,705,1176,1785,1937,2219,2503,2865,3921,3945,
0,11,277,306,332,968,1477,1624,2048,2494,2905,3128,4184,4208,
134,205,287,326,991,1067,1728,1993,2071,2301,3151,3189,4207,4231,
23,137,201,281,375,569,1347,1361,1373,2336,2441,2937,3497,3521,
110,194,211,258,298,504,1274,1331,2159,2327,2354,2784,3410,3434,
128,202,263,485,655,926,1104,1565,1798,2645,2727,3188,3701,3725,
7,59,92,152,243,750,1087,1428,1676,2167,2258,3037,3247,4302,
39,63,106,270,386,515,1367,1595,1969,2488,2649,2675,3731,3755,
137,164,200,224,306,394,1174,1244,2138,2324,2361,2551,3380,3404,
36,47,76,580,589,1014,1309,1533,2094,2249,2825,3174,4230,4254,
90,142,170,198,213,423,1170,1172,1207,2250,2973,3218,3306,3330,
154,208,222,498,667,831,1133,1747,1770,2340,2827,2845,3883,3907,
203,235,277,535,605,1022,1685,1897,1955,2211,2765,2841,3821,3845,
7,172,263,459,781,938,1195,2007,2018,2437,2685,3098,4154,4178,
46,234,294,321,342,905,1318,1843,1985,2430,3065,3215,4121,4145,
164,166,191,274,337,442,1210,1449,1522,2602,2870,2923,3658,3682,
4,142,206,286,380,574,1352,1366,1378,2341,2446,2942,3502,3526,
23,105,177,326,755,1056,1420,1723,1835,2396,2915,3217,3971,3995,
246,344,355,607,693,1055,1726,1773,1818,2689,2853,3094,3909,3933,
9,174,241,461,783,940,1197,2009,2020,2439,2687,3100,4156,4180,
11,176,243,463,785,942,1199,2011,2022,2441,2665,3102,4158,4182,
38,69,87,214,427,771,1085,1687,1851,2879,2931,3067,3987,4011,
154,156,181,264,351,432,1200,1463,1512,2592,2860,2913,3648,3672,
30,51,97,151,217,700,1297,1381,2111,2377,2610,2672,3433,3457,
104,205,212,252,292,522,1292,1325,2153,2321,2372,2802,3428,3452,
6,69,294,305,332,753,1255,1374,1833,2161,2454,2496,3510,3534,
138,165,201,225,307,395,1175,1245,2139,2325,2362,2552,3381,3405,
134,161,197,221,303,391,1171,1241,2159,2321,2358,2548,3377,3401,
14,135,283,301,433,717,1188,1797,1925,2231,2515,2877,3933,3957,
247,345,356,608,694,1032,1727,1774,1819,2690,2854,3095,3910,3934,
26,48,111,278,992,1045,1747,1788,2125,2769,2777,3205,4261,4285,
6,171,262,458,780,937,1194,2006,2017,2436,2684,3097,4153,4177,
119,191,240,362,449,634,1442,1648,2085,2467,2522,3018,3578,3602,
41,229,289,316,337,900,1313,1838,1980,2425,3060,3210,4116,4140,
143,193,254,500,670,917,1119,1580,1789,2660,2718,3179,3716,3740,
1,122,159,565,573,885,1334,1538,1653,2550,2625,2733,3789,3813,
47,69,108,275,989,1042,1744,1785,2122,2766,2774,3202,4258,4282,
29,42,82,586,595,1020,1315,1515,2100,2255,2831,3180,4236,4260,
25,48,55,173,729,980,1135,1247,2056,2178,2215,2747,3271,3295,
27,239,299,326,347,910,1299,1824,1990,2435,3070,3196,4126,4150,
15,129,193,273,367,561,1353,1363,1389,2328,2433,2929,3489,3513,
29,92,188,223,959,976,1109,1489,1980,2189,2722,3113,3245,3269,
144,146,171,278,341,446,1214,1453,1526,2606,2874,2927,3662,3686,
33,97,226,253,292,314,1333,1514,1877,2388,2413,2421,3469,3493,
31,219,303,330,351,890,1303,1828,1970,2439,3050,3200,4106,4130,
98,170,243,365,452,637,1445,1651,2064,2470,2525,3021,3581,3605,
123,133,140,226,742,778,1203,1759,1870,2276,2283,3147,3339,3363,
185,240,355,520,799,922,1554,2002,2122,3001,3082,3129,4138,4162,
87,110,307,319,349,530,1240,1429,1494,2509,2542,2799,3565,3589,
18,139,287,305,437,697,1192,1777,1929,2211,2519,2857,3913,3937,
124,131,138,217,733,769,1218,1774,1861,2267,2298,3162,3354,3378,
9,55,104,200,219,549,1629,1950,2023,2361,2709,2902,3765,3789,
2,140,204,284,378,572,1350,1364,1376,2339,2444,2940,3500,3524,
127,198,280,319,984,1060,1745,2010,2064,2294,3144,3182,4200,4224,
7,70,295,306,333,754,1256,1375,1834,2162,2455,2497,3511,3535,
89,148,151,226,395,854,1475,2030,2055,2204,2555,2757,3611,3635,
187,242,357,522,801,924,1556,2004,2124,3003,3084,3131,4140,4164,
188,219,326,343,460,809,1136,1268,1589,2348,2606,2961,3404,3428,
29,50,96,150,216,699,1296,1380,2110,2376,2609,2671,3432,3456,
33,72,168,227,939,980,1113,1493,1984,2193,2726,3117,3249,3273,
7,128,165,555,571,867,1340,1544,1635,2556,2631,2715,3771,3795,
110,255,274,316,334,1003,1284,1396,1645,2476,2589,2652,3532,3556,
85,108,305,317,347,528,1238,1427,1492,2507,2540,2797,3563,3587,
63,96,251,277,697,871,1100,1112,1176,2256,2404,2571,3312,3336,
98,243,286,322,328,991,1272,1408,1633,2488,2577,2640,3544,3568,
125,135,142,228,720,780,1205,1761,1848,2278,2285,3149,3341,3365,
10,23,276,305,331,967,1476,1623,2047,2493,2904,3127,4183,4207,
94,122,174,193,202,427,1152,1174,1211,2254,2953,3222,3310,3334,
190,221,328,345,462,811,1138,1270,1591,2350,2608,2963,3406,3430,
71,180,305,819,825,898,1406,1486,1905,2527,2618,2985,4041,4065,
17,63,112,208,227,533,1613,1958,2031,2369,2693,2886,3749,3773,
32,43,72,576,585,1010,1305,1529,2090,2245,2821,3170,4226,4250,
75,158,161,236,405,840,1485,2016,2041,2190,2565,2743,3621,3645,
76,121,272,351,645,852,1285,1932,2071,2705,2942,3012,4068,4092,
241,339,350,602,688,1050,1721,1768,1813,2708,2848,3089,3904,3928,
159,213,227,503,648,836,1138,1728,1775,2345,2808,2850,3864,3888,
30,177,293,361,1048,1078,1462,1802,2158,2240,3151,3238,4294,4318,
251,348,357,812,911,1010,1263,1576,1892,2288,2972,3129,4028,4052,
258,340,355,795,894,1017,1270,1583,1875,2295,2955,3136,4011,4035,
24,35,88,577,592,1026,1297,1521,2106,2237,2813,3186,4242,4266,
27,51,118,282,398,527,1355,1607,1981,2476,2661,2687,3743,3767,
212,220,286,544,614,1031,1694,1906,1964,2220,2774,2850,3830,3854,
83,121,157,313,683,881,1606,1917,1961,2817,2983,3041,4097,4121,
80,163,166,217,386,845,1466,2021,2046,2195,2546,2748,3602,3626,
65,98,253,279,699,873,1102,1114,1178,2258,2406,2573,3314,3338,
162,164,189,272,359,440,1208,1447,1520,2600,2868,2921,3656,3680,
70,103,258,284,704,878,1083,1119,1183,2263,2411,2578,3319,3343,
91,150,153,228,397,856,1477,2032,2057,2206,2557,2759,3613,3637,
31,178,294,362,1049,1079,1463,1803,2159,2241,3152,3239,4295,4319,
23,191,341,347,613,630,1409,1625,1710,2790,2902,3073,3846,3870,
45,52,94,197,410,778,1092,1694,1858,2862,2938,3050,3994,4018,
27,50,57,175,731,982,1137,1225,2058,2180,2217,2749,3273,3297,
67,84,85,427,691,953,1507,1679,2127,2456,2587,3105,3643,3667,
18,139,152,558,566,878,1327,1555,1646,2567,2618,2726,3782,3806,
249,347,358,610,672,1034,1705,1752,1821,2692,2832,3073,3888,3912,
25,88,184,219,955,972,1105,1509,1976,2185,2718,3109,3241,3265,
83,135,187,206,215,416,1163,1165,1200,2243,2966,3235,3299,3323,
129,136,143,222,738,774,1223,1755,1866,2272,2303,3167,3359,3383,
101,173,246,368,455,640,1448,1654,2067,2449,2528,3000,3584,3608,
11,63,72,156,247,754,1091,1432,1656,2171,2262,3041,3251,4306,
94,139,266,345,639,846,1279,1926,2065,2699,2936,3006,4062,4086,
6,17,283,288,314,974,1483,1630,2054,2476,2911,3134,4190,4214,
180,235,318,359,476,801,1128,1260,1605,2340,2598,2953,3396,3420,
146,200,238,490,659,823,1149,1739,1762,2332,2819,2837,3875,3899,
92,151,154,229,398,857,1478,2033,2058,2207,2558,2736,3614,3638,
60,77,78,420,684,946,1500,1672,2120,2449,2580,3098,3636,3660,
255,337,352,792,891,1014,1267,1580,1872,2292,2952,3133,4008,4032,
19,140,264,306,438,698,1193,1778,1930,2212,2496,2858,3914,3938,
117,194,201,241,305,511,1281,1338,2142,2310,2361,2791,3417,3441,
36,60,103,267,407,512,1364,1592,1990,2485,2646,2672,3728,3752,
28,39,92,581,596,1030,1301,1525,2110,2241,2817,3190,4246,4270,
153,207,221,497,666,830,1132,1746,1769,2339,2826,2844,3882,3906,
86,124,160,316,686,884,1585,1896,1964,2820,2986,3044,4100,4124,
260,345,358,621,683,1045,1716,1763,1808,2703,2843,3084,3899,3923,
45,84,180,239,951,968,1125,1505,1972,2205,2714,3105,3261,3285,
92,137,264,343,637,844,1277,1924,2087,2697,2934,3004,4060,4084,
4,125,162,552,568,864,1337,1541,1632,2553,2628,2712,3768,3792,
7,121,209,265,383,553,1345,1355,1381,2344,2425,2945,3481,3505,
257,339,354,794,893,1016,1269,1582,1874,2294,2954,3135,4010,4034,
60,117,248,274,718,868,1097,1109,1197,2277,2401,2568,3333,3357,
26,39,79,583,592,1017,1312,1512,2097,2252,2828,3177,4233,4257,
32,95,191,226,938,979,1112,1492,1983,2192,2725,3116,3248,3272,
18,186,336,342,608,625,1404,1620,1705,2785,2897,3092,3841,3865,
100,201,208,248,288,518,1288,1321,2149,2317,2368,2798,3424,3448,
89,144,159,246,492,723,1562,1680,1803,2192,2883,3028,3939,3963,
204,236,278,536,606,1023,1686,1898,1956,2212,2766,2842,3822,3846,
39,227,311,314,359,898,1311,1836,1978,2447,3058,3208,4114,4138,
44,232,292,319,340,903,1316,1841,1983,2428,3063,3213,4119,4143,
92,120,172,200,215,425,1172,1174,1209,2252,2975,3220,3308,3332,
17,99,171,320,749,1074,1438,1717,1829,2390,2909,3235,3965,3989,
149,203,217,493,662,826,1128,1742,1765,2335,2822,2840,3878,3902,
3,141,205,285,379,573,1351,1365,1377,2340,2445,2941,3501,3525,
43,50,92,195,408,776,1090,1692,1856,2860,2936,3048,3992,4016,
15,237,272,576,661,914,1656,1894,1935,2736,2997,3209,3792,3816,
191,222,329,346,463,812,1139,1271,1592,2351,2609,2964,3407,3431,
150,204,218,494,663,827,1129,1743,1766,2336,2823,2841,3879,3903,
74,136,148,328,674,872,1597,1908,1952,2808,2998,3032,4088,4112,
76,99,296,332,338,543,1229,1418,1507,2498,2531,2788,3554,3578,
210,218,284,542,612,1029,1692,1904,1962,2218,2772,2848,3828,3852,
30,43,83,587,596,1021,1316,1516,2101,2232,2808,3181,4237,4261,
37,68,86,213,426,770,1084,1686,1850,2878,2930,3066,3986,4010,
36,58,97,264,1002,1055,1733,1798,2135,2763,2779,3215,4271,4295,
131,158,194,218,300,388,1168,1238,2156,2318,2355,2545,3374,3398,
79,124,275,354,624,855,1288,1935,2074,2708,2945,3015,4071,4095,
11,57,106,202,221,551,1631,1952,2025,2363,2711,2880,3767,3791,
21,189,339,345,611,628,1407,1623,1708,2788,2900,3095,3844,3868,
9,130,278,296,452,712,1183,1792,1920,2226,2510,2872,3928,3952,
38,60,99,266,1004,1033,1735,1776,2113,2765,2781,3193,4249,4273,
122,129,136,239,731,791,1216,1772,1859,2265,2296,3160,3352,3376,
120,127,137,230,722,782,1207,1763,1850,2256,2287,3151,3343,3367,
182,237,320,337,478,803,1130,1262,1607,2342,2600,2955,3398,3422,
34,98,227,254,293,315,1334,1515,1878,2389,2414,2422,3470,3494,
169,224,331,348,465,814,1141,1249,1594,2329,2611,2966,3385,3409,
128,135,142,221,737,773,1222,1754,1865,2271,2302,3166,3358,3382,
81,164,167,218,387,846,1467,2022,2047,2196,2547,2749,3603,3627,
20,141,265,307,439,699,1194,1779,1931,2213,2497,2859,3915,3939,
43,65,104,271,985,1038,1740,1781,2118,2762,2770,3198,4254,4278,
54,72,95,414,678,940,1494,1666,2114,2467,2574,3116,3630,3654,
32,63,81,208,421,789,1103,1681,1869,2873,2949,3061,4005,4029,
22,187,254,474,772,953,1186,1998,2033,2428,2676,3113,4169,4193,
78,101,298,334,340,545,1231,1420,1509,2500,2533,2790,3556,3580,
3,124,272,290,446,706,1177,1786,1938,2220,2504,2866,3922,3946,
21,142,155,561,569,881,1330,1558,1649,2546,2621,2729,3785,3809,
40,63,70,188,720,971,1150,1238,2047,2169,2230,2738,3286,3310,
95,150,165,252,498,729,1568,1686,1809,2198,2889,3034,3945,3969,
14,135,148,554,562,874,1323,1551,1642,2563,2638,2722,3778,3802,
16,137,285,303,435,719,1190,1799,1927,2209,2517,2879,3935,3959,
28,59,77,204,417,785,1099,1701,1865,2869,2945,3057,4001,4025,
144,198,236,488,657,821,1147,1737,1760,2330,2817,2835,3873,3897,
11,132,145,559,575,871,1320,1548,1639,2560,2635,2719,3775,3799,
15,54,290,303,317,762,1264,1383,1842,2170,2463,2505,3519,3543,
16,238,273,577,662,915,1657,1895,1936,2737,2998,3210,3793,3817,
117,189,262,360,447,632,1440,1646,2083,2465,2520,3016,3576,3600,
161,163,188,271,358,439,1207,1446,1519,2599,2867,2920,3655,3679,
27,174,290,382,1045,1075,1459,1823,2155,2237,3148,3235,4291,4315,
135,206,264,327,992,1068,1729,1994,2072,2302,3152,3190,4208,4232,
30,118,223,250,289,335,1330,1535,1874,2385,2410,2418,3466,3490,
4,110,182,331,760,1061,1425,1704,1840,2377,2920,3222,3976,4000,
123,197,258,480,650,921,1123,1560,1793,2640,2722,3183,3696,3720,
72,151,166,253,499,730,1569,1687,1810,2199,2890,3035,3946,3970,
17,138,286,304,436,696,1191,1776,1928,2210,2518,2856,3912,3936,
36,183,299,367,1054,1060,1444,1808,2140,2246,3157,3220,4276,4300,
77,122,273,352,646,853,1286,1933,2072,2706,2943,3013,4069,4093,
163,193,231,483,652,816,1142,1732,1755,2349,2812,2854,3868,3892,
215,223,265,547,617,1010,1697,1909,1967,2223,2777,2853,3833,3857,
33,64,82,209,422,790,1080,1682,1870,2874,2950,3062,4006,4030,
111,183,256,378,441,626,1458,1640,2077,2459,2538,3010,3594,3618,
12,118,190,315,744,1069,1433,1712,1824,2385,2904,3230,3960,3984,
39,70,88,215,428,772,1086,1688,1852,2856,2932,3068,3988,4012,
34,55,101,155,221,704,1301,1385,2091,2381,2614,2676,3437,3461,
66,99,254,280,700,874,1103,1115,1179,2259,2407,2574,3315,3339,
171,250,341,506,809,932,1540,2012,2132,3011,3092,3139,4148,4172,
78,140,152,332,678,876,1601,1912,1956,2812,2978,3036,4092,4116,
116,188,261,383,446,631,1463,1645,2082,2464,2543,3015,3599,3623,
72,124,176,195,204,429,1152,1154,1213,2232,2955,3224,3288,3312,
31,54,61,179,735,962,1141,1229,2062,2160,2221,2753,3277,3301,
22,220,279,583,668,921,1663,1877,1942,2743,2980,3192,3799,3823,
240,338,349,601,687,1049,1720,1767,1812,2707,2847,3088,3903,3927,
147,201,239,491,660,824,1150,1740,1763,2333,2820,2838,3876,3900,
109,181,254,376,439,624,1456,1638,2075,2457,2536,3008,3592,3616,
33,54,100,154,220,703,1300,1384,2090,2380,2613,2675,3436,3460,
75,127,179,198,207,408,1155,1157,1216,2235,2958,3227,3291,3315,
61,118,249,275,719,869,1098,1110,1198,2278,2402,2569,3334,3358,
156,210,224,500,669,833,1135,1749,1772,2342,2829,2847,3885,3909,
83,145,166,220,389,848,1469,2024,2049,2198,2549,2751,3605,3629,
8,114,186,335,764,1065,1429,1708,1844,2381,2924,3226,3980,4004,
88,147,150,225,394,853,1474,2029,2054,2203,2554,2756,3610,3634,
30,102,307,320,474,860,1554,1860,2098,2315,2634,3051,3690,3714,
35,57,96,287,1001,1054,1732,1797,2134,2762,2778,3214,4270,4294,
86,156,165,243,489,720,1583,1701,1800,2189,2880,3025,3936,3960,
158,212,226,502,671,835,1137,1751,1774,2344,2831,2849,3887,3911,
58,115,246,272,716,866,1095,1107,1195,2275,2423,2590,3331,3355,
186,241,356,521,800,923,1555,2003,2123,3002,3083,3130,4139,4163,
40,62,101,268,1006,1035,1737,1778,2115,2767,2783,3195,4251,4275,
123,194,276,315,1004,1056,1741,2006,2084,2290,3164,3178,4220,4244,
120,127,134,237,729,789,1214,1770,1857,2263,2294,3158,3350,3374,
1,12,278,307,333,969,1478,1625,2049,2495,2906,3129,4185,4209,
86,138,190,194,209,419,1166,1168,1203,2246,2969,3238,3302,3326,
25,70,116,146,236,719,1316,1376,2106,2396,2605,2667,3452,3476,
122,193,275,314,1003,1079,1740,2005,2083,2289,3163,3177,4219,4243,
62,119,250,276,696,870,1099,1111,1199,2279,2403,2570,3335,3359,
3,16,269,298,324,960,1469,1616,2040,2486,2921,3120,4176,4200,
85,130,281,336,630,861,1294,1941,2080,2690,2951,3021,4077,4101,
107,208,215,255,295,525,1295,1328,2156,2324,2375,2805,3431,3455,
5,57,90,150,241,748,1085,1426,1674,2165,2256,3035,3245,4300,
56,113,244,270,714,864,1093,1105,1193,2273,2421,2588,3329,3353,
247,344,353,808,907,1030,1259,1572,1888,2284,2968,3125,4024,4048,
86,145,148,223,392,851,1472,2027,2052,2201,2552,2754,3608,3632,
262,336,347,623,685,1047,1718,1765,1810,2705,2845,3086,3901,3925,
243,341,352,604,690,1052,1723,1770,1815,2710,2850,3091,3906,3930,
76,128,180,199,208,409,1156,1158,1217,2236,2959,3228,3292,3316,
135,162,198,222,304,392,1172,1242,2136,2322,2359,2549,3378,3402,
71,104,259,285,705,879,1084,1120,1184,2264,2412,2579,3320,3344,
79,141,153,333,679,877,1602,1913,1957,2813,2979,3037,4093,4117,
44,191,307,375,1038,1068,1452,1816,2148,2254,3165,3228,4284,4308,
3,124,161,567,575,887,1336,1540,1655,2552,2627,2735,3791,3815,
54,187,288,826,832,905,1413,1469,1912,2534,2625,2992,4048,4072,
25,71,110,277,991,1044,1746,1787,2124,2768,2776,3204,4260,4284,
149,151,176,283,346,451,1219,1458,1531,2611,2879,2908,3667,3691,
47,119,300,313,467,853,1547,1853,2091,2308,2627,3068,3683,3707,
200,232,274,532,602,1019,1682,1918,1952,2208,2762,2838,3818,3842,
87,132,283,338,632,863,1272,1943,2082,2692,2929,3023,4079,4103,
16,55,291,304,318,763,1265,1384,1843,2171,2464,2506,3520,3544,
141,212,270,333,998,1074,1735,2000,2078,2284,3158,3172,4214,4238,
6,19,272,301,327,963,1472,1619,2043,2489,2924,3123,4179,4203,
199,231,273,531,601,1018,1681,1917,1951,2231,2761,2837,3817,3841,
77,139,151,331,677,875,1600,1911,1955,2811,2977,3035,4091,4115,
166,196,234,486,655,819,1145,1735,1758,2328,2815,2833,3871,3895,
170,225,332,349,466,815,1142,1250,1595,2330,2612,2967,3386,3410,
34,222,306,333,354,893,1306,1831,1973,2442,3053,3203,4109,4133,
81,133,185,204,213,414,1161,1163,1222,2241,2964,3233,3297,3321,
13,52,288,301,315,760,1262,1381,1840,2168,2461,2503,3517,3541,
14,236,271,599,660,913,1679,1893,1934,2759,2996,3208,3815,3839,
59,168,293,831,837,910,1394,1474,1917,2539,2630,2997,4053,4077,
32,96,225,252,291,313,1332,1513,1876,2387,2412,2420,3468,3492,
148,202,216,492,661,825,1151,1741,1764,2334,2821,2839,3877,3901,
28,116,221,248,311,333,1328,1533,1872,2383,2408,2416,3464,3488,
12,177,244,464,786,943,1176,2012,2023,2442,2666,3103,4159,4183,
37,59,98,265,1003,1032,1734,1799,2112,2764,2780,3192,4248,4272,
74,143,270,349,643,850,1283,1930,2069,2703,2940,3010,4066,4090,
0,70,119,215,234,540,1620,1965,2038,2352,2700,2893,3756,3780,
50,91,92,410,674,936,1490,1662,2134,2463,2570,3112,3626,3650,
85,144,147,222,391,850,1471,2026,2051,2200,2551,2753,3607,3631,
33,180,296,364,1051,1057,1441,1805,2137,2243,3154,3217,4273,4297,
142,192,253,499,669,916,1118,1579,1788,2659,2717,3178,3715,3739,
7,53,102,198,217,547,1627,1948,2021,2359,2707,2900,3763,3787,
30,52,115,282,996,1049,1751,1792,2129,2773,2781,3209,4265,4289,
78,161,164,239,384,843,1464,2019,2044,2193,2544,2746,3600,3624,
24,87,183,218,954,971,1104,1508,1975,2184,2717,3108,3240,3264,
18,64,113,209,228,534,1614,1959,2032,2370,2694,2887,3750,3774,
22,143,267,309,441,701,1196,1781,1933,2215,2499,2861,3917,3941,
28,175,291,383,1046,1076,1460,1800,2156,2238,3149,3236,4292,4316,
30,53,60,178,734,961,1140,1228,2061,2183,2220,2752,3276,3300,
21,186,253,473,771,952,1185,1997,2032,2427,2675,3112,4168,4192,
82,127,278,357,627,858,1291,1938,2077,2711,2948,3018,4074,4098,
42,66,109,273,389,518,1346,1598,1972,2491,2652,2678,3734,3758,
25,36,89,578,593,1027,1298,1522,2107,2238,2814,3187,4243,4267,
23,120,268,310,442,702,1197,1782,1934,2216,2500,2862,3918,3942,
16,68,77,161,252,759,1096,1437,1661,2176,2267,3046,3256,4311,
254,339,352,615,677,1039,1710,1757,1802,2697,2837,3078,3893,3917,
128,199,281,320,985,1061,1746,2011,2065,2295,3145,3183,4201,4225,
12,133,146,552,560,872,1321,1549,1640,2561,2636,2720,3776,3800,
37,60,67,185,741,968,1147,1235,2044,2166,2227,2759,3283,3307,
145,147,172,279,342,447,1215,1454,1527,2607,2875,2904,3663,3687,
32,55,62,180,736,963,1142,1230,2063,2161,2222,2754,3278,3302,
26,238,298,325,346,909,1298,1847,1989,2434,3069,3195,4125,4149,
11,22,264,293,319,979,1464,1611,2059,2481,2916,3139,4195,4219,
28,41,81,585,594,1019,1314,1514,2099,2254,2830,3179,4235,4259,
172,251,342,507,810,933,1541,2013,2133,3012,3093,3140,4149,4173,
87,146,149,224,393,852,1473,2028,2053,2202,2553,2755,3609,3633,
167,197,235,487,656,820,1146,1736,1759,2329,2816,2834,3872,3896,
48,89,90,408,672,958,1488,1660,2132,2461,2568,3110,3624,3648,
25,97,302,315,469,855,1549,1855,2093,2310,2629,3070,3685,3709,
28,49,119,149,239,698,1319,1379,2109,2399,2608,2670,3455,3479,
31,62,80,207,420,788,1102,1680,1868,2872,2948,3060,4004,4028,
8,173,240,460,782,939,1196,2008,2019,2438,2686,3099,4155,4179,
51,108,263,265,709,883,1088,1124,1188,2268,2416,2583,3324,3348,
40,79,175,234,946,963,1120,1500,1991,2200,2733,3100,3256,3280,
81,126,277,356,626,857,1290,1937,2076,2710,2947,3017,4073,4097,
9,22,275,304,330,966,1475,1622,2046,2492,2927,3126,4182,4206,
17,56,292,305,319,764,1266,1385,1844,2172,2465,2507,3521,3545,
85,155,164,242,488,743,1582,1700,1823,2188,2903,3024,3959,3983,
28,51,58,176,732,983,1138,1226,2059,2181,2218,2750,3274,3298,
107,179,252,374,437,646,1454,1636,2073,2455,2534,3006,3590,3614,
47,235,295,322,343,906,1319,1844,1986,2431,3066,3192,4122,4146,
25,237,297,324,345,908,1297,1846,1988,2433,3068,3194,4124,4148,
208,216,282,540,610,1027,1690,1902,1960,2216,2770,2846,3826,3850,
11,132,280,298,454,714,1185,1794,1922,2228,2512,2874,3930,3954,
39,62,69,187,743,970,1149,1237,2046,2168,2229,2737,3285,3309,
82,105,302,314,344,549,1235,1424,1489,2504,2537,2794,3560,3584,
45,109,238,241,304,326,1321,1526,1889,2376,2401,2409,3457,3481,
76,159,162,237,406,841,1486,2017,2042,2191,2566,2744,3622,3646,
141,144,204,228,310,398,1154,1224,2142,2304,2365,2555,3360,3384,
14,128,192,272,366,560,1352,1362,1388,2351,2432,2928,3488,3512,
31,44,84,588,597,1022,1317,1517,2102,2233,2809,3182,4238,4262,
34,45,74,578,587,1012,1307,1531,2092,2247,2823,3172,4228,4252,
190,245,336,525,804,927,1559,2007,2127,3006,3087,3134,4143,4167,
252,349,358,813,888,1011,1264,1577,1893,2289,2973,3130,4029,4053,
83,153,162,240,486,741,1580,1698,1821,2186,2901,3046,3957,3981,
138,209,267,330,995,1071,1732,1997,2075,2281,3155,3169,4211,4235,
38,185,301,369,1032,1062,1446,1810,2142,2248,3159,3222,4278,4302,
44,108,237,240,303,325,1320,1525,1888,2399,2400,2408,3456,3480,
42,64,103,270,984,1037,1739,1780,2117,2761,2769,3197,4253,4277,
19,101,173,322,751,1076,1416,1719,1831,2392,2911,3237,3967,3991,
12,58,107,203,222,528,1608,1953,2026,2364,2688,2881,3744,3768,
36,57,103,157,223,706,1303,1387,2093,2383,2592,2678,3439,3463,
189,220,327,344,461,810,1137,1269,1590,2349,2607,2962,3405,3429,
6,112,184,333,762,1063,1427,1706,1842,2379,2922,3224,3978,4002,
88,111,308,320,350,531,1241,1430,1495,2510,2543,2800,3566,3590,
52,109,240,266,710,884,1089,1125,1189,2269,2417,2584,3325,3349,
3,171,345,351,617,634,1413,1629,1714,2794,2882,3077,3850,3874,
123,130,137,216,732,768,1217,1773,1860,2266,2297,3161,3353,3377,
36,100,229,256,295,317,1336,1517,1880,2391,2400,2416,3472,3496,
12,51,300,311,314,759,1261,1380,1839,2167,2460,2502,3516,3540,
198,230,272,530,600,1017,1680,1916,1950,2230,2760,2836,3816,3840,
105,206,213,253,293,523,1293,1326,2154,2322,2373,2803,3429,3453,
46,169,309,377,1040,1070,1454,1818,2150,2232,3167,3230,4286,4310,
94,117,290,326,356,537,1247,1436,1501,2516,2525,2806,3572,3596,
20,48,81,165,256,763,1100,1417,1665,2180,2271,3026,3260,4315,
8,21,274,303,329,965,1474,1621,2045,2491,2926,3125,4181,4205,
37,225,309,312,357,896,1309,1834,1976,2445,3056,3206,4112,4136,
19,65,114,210,229,535,1615,1960,2033,2371,2695,2888,3751,3775,
79,149,158,260,482,737,1576,1694,1817,2206,2897,3042,3953,3977,
82,144,165,219,388,847,1468,2023,2048,2197,2548,2750,3604,3628,
92,130,166,322,692,866,1591,1902,1946,2826,2992,3026,4082,4106,
93,138,265,344,638,845,1278,1925,2064,2698,2935,3005,4061,4085,
34,73,169,228,940,981,1114,1494,1985,2194,2727,3118,3250,3274,
47,111,216,243,306,328,1323,1528,1891,2378,2403,2411,3459,3483,
70,87,88,430,694,956,1510,1658,2130,2459,2590,3108,3646,3670,
172,227,334,351,468,793,1144,1252,1597,2332,2614,2969,3388,3412,
261,343,358,798,897,1020,1249,1562,1878,2298,2958,3139,4014,4038,
144,166,169,276,339,444,1212,1451,1524,2604,2872,2925,3660,3684,
175,230,313,354,471,796,1147,1255,1600,2335,2593,2972,3391,3415,
140,211,269,332,997,1073,1734,1999,2077,2283,3157,3171,4213,4237,
152,154,179,286,349,454,1222,1461,1534,2614,2858,2911,3670,3694,
244,341,350,805,904,1027,1256,1569,1885,2281,2965,3122,4021,4045,
119,240,283,319,325,988,1293,1405,1654,2485,2574,2661,3541,3565,
68,101,256,282,702,876,1081,1117,1181,2261,2409,2576,3317,3341,
29,52,59,177,733,960,1139,1227,2060,2182,2219,2751,3275,3299,
136,163,199,223,305,393,1173,1243,2137,2323,2360,2550,3379,3403,
95,118,291,327,357,538,1224,1437,1502,2517,2526,2807,3573,3597,
39,78,174,233,945,962,1119,1499,1990,2199,2732,3099,3255,3279,
19,217,276,580,665,918,1660,1874,1939,2740,2977,3213,3796,3820,
126,133,143,236,728,788,1213,1769,1856,2262,2293,3157,3349,3373,
111,256,275,317,335,1004,1285,1397,1646,2477,2590,2653,3533,3557,
30,54,97,285,401,506,1358,1586,1984,2479,2640,2666,3722,3746,
37,58,104,158,224,707,1304,1388,2094,2384,2593,2679,3440,3464,
49,182,307,821,827,900,1408,1464,1907,2529,2620,2987,4043,4067,
64,81,82,424,688,950,1504,1676,2124,2453,2584,3102,3640,3664,
38,226,310,313,358,897,1310,1835,1977,2446,3057,3207,4113,4137,
170,249,340,505,808,931,1539,2011,2131,3010,3091,3138,4147,4171,
126,153,213,237,295,407,1163,1233,2151,2313,2374,2564,3369,3393,
80,142,154,334,680,878,1603,1914,1958,2814,2980,3038,4094,4118,
20,188,338,344,610,627,1406,1622,1707,2787,2899,3094,3843,3867,
171,226,333,350,467,792,1143,1251,1596,2331,2613,2968,3387,3411,
2,108,180,329,758,1059,1423,1726,1838,2399,2918,3220,3974,3998,
6,228,287,591,652,929,1671,1885,1926,2751,2988,3200,3807,3831,
0,138,202,282,376,570,1348,1362,1374,2337,2442,2938,3498,3522,
145,167,170,277,340,445,1213,1452,1525,2605,2873,2926,3661,3685,
23,188,255,475,773,954,1187,1999,2034,2429,2677,3114,4170,4194,
168,247,338,527,806,929,1537,2009,2129,3008,3089,3136,4145,4169,
47,54,72,199,412,780,1094,1696,1860,2864,2940,3052,3996,4020,
20,59,295,308,322,767,1269,1388,1847,2175,2468,2510,3524,3548,
136,210,247,493,663,934,1112,1573,1782,2653,2735,3172,3709,3733,
25,38,78,582,591,1016,1311,1535,2096,2251,2827,3176,4232,4256,
101,202,209,249,289,519,1289,1322,2150,2318,2369,2799,3425,3449,
29,176,292,360,1047,1077,1461,1801,2157,2239,3150,3237,4293,4317,
100,245,264,324,330,993,1274,1410,1635,2490,2579,2642,3546,3570,
9,177,351,357,623,640,1395,1611,1720,2800,2888,3083,3856,3880,
88,126,162,318,688,886,1587,1898,1966,2822,2988,3046,4102,4126,
5,227,286,590,651,928,1670,1884,1925,2750,2987,3199,3806,3830,
89,134,285,340,634,841,1274,1921,2084,2694,2931,3001,4057,4081,
242,339,348,803,902,1025,1254,1567,1883,2303,2963,3120,4019,4043,
2,13,279,308,334,970,1479,1626,2050,2472,2907,3130,4186,4210,
52,93,94,412,676,938,1492,1664,2112,2465,2572,3114,3628,3652,
155,209,223,499,668,832,1134,1748,1771,2341,2828,2846,3884,3908,
143,214,272,335,1000,1076,1737,2002,2080,2286,3160,3174,4216,4240,
254,336,351,815,890,1013,1266,1579,1895,2291,2975,3132,4031,4055,
132,159,195,219,301,389,1169,1239,2157,2319,2356,2546,3375,3399,
33,56,63,181,737,964,1143,1231,2040,2162,2223,2755,3279,3303,
75,120,271,350,644,851,1284,1931,2070,2704,2941,3011,4067,4091,
17,239,274,578,663,916,1658,1872,1937,2738,2999,3211,3794,3818,
106,207,214,254,294,524,1294,1327,2155,2323,2374,2804,3430,3454,
33,44,73,577,586,1011,1306,1530,2091,2246,2822,3171,4227,4251,
43,231,291,318,339,902,1315,1840,1982,2427,3062,3212,4118,4142,
17,69,78,162,253,760,1097,1438,1662,2177,2268,3047,3257,4312,
8,71,296,307,334,755,1257,1376,1835,2163,2456,2498,3512,3536,
42,63,109,163,229,712,1309,1369,2099,2389,2598,2684,3445,3469,
55,112,243,269,713,887,1092,1104,1192,2272,2420,2587,3328,3352,
40,228,288,315,336,899,1312,1837,1979,2424,3059,3209,4115,4139,
86,109,306,318,348,529,1239,1428,1493,2508,2541,2798,3564,3588,
73,135,147,327,673,871,1596,1907,1951,2831,2997,3031,4087,4111,
32,220,304,331,352,891,1304,1829,1971,2440,3051,3201,4107,4131,
177,256,347,512,815,914,1546,1994,2114,3017,3074,3121,4130,4154,
50,107,262,264,708,882,1087,1123,1187,2267,2415,2582,3323,3347,
31,94,190,225,937,978,1111,1491,1982,2191,2724,3115,3247,3271,
256,341,354,617,679,1041,1712,1759,1804,2699,2839,3080,3895,3919,
214,222,264,546,616,1009,1696,1908,1966,2222,2776,2852,3832,3856,
125,132,142,235,727,787,1212,1768,1855,2261,2292,3156,3348,3372,
79,131,183,202,211,412,1159,1161,1220,2239,2962,3231,3295,3319,
35,99,228,255,294,316,1335,1516,1879,2390,2415,2423,3471,3495,
30,93,189,224,936,977,1110,1490,1981,2190,2723,3114,3246,3270,
82,152,161,263,485,740,1579,1697,1820,2185,2900,3045,3956,3980,
12,133,281,299,455,715,1186,1795,1923,2229,2513,2875,3931,3955,
6,52,101,197,216,546,1626,1947,2020,2358,2706,2899,3762,3786,
97,242,285,321,327,990,1295,1407,1632,2487,2576,2663,3543,3567,
241,338,347,802,901,1024,1253,1566,1882,2302,2962,3143,4018,4042,
262,344,359,799,898,1021,1250,1563,1879,2299,2959,3140,4015,4039,
9,20,286,291,317,977,1486,1609,2057,2479,2914,3137,4193,4217,
10,131,279,297,453,713,1184,1793,1921,2227,2511,2873,3929,3953,
92,147,162,249,495,726,1565,1683,1806,2195,2886,3031,3942,3966,
98,199,206,246,310,516,1286,1343,2147,2315,2366,2796,3422,3446,
6,127,164,554,570,866,1339,1543,1634,2555,2630,2714,3770,3794,
12,64,73,157,248,755,1092,1433,1657,2172,2263,3042,3252,4307,
8,129,166,556,572,868,1341,1545,1636,2557,2632,2716,3772,3796,
109,254,273,315,333,1002,1283,1395,1644,2475,2588,2651,3531,3555,
5,18,271,300,326,962,1471,1618,2042,2488,2923,3122,4178,4202,
24,236,296,323,344,907,1296,1845,1987,2432,3067,3193,4123,4147,
35,223,307,334,355,894,1307,1832,1974,2443,3054,3204,4110,4134,
9,48,297,308,335,756,1258,1377,1836,2164,2457,2499,3513,3537,
81,104,301,313,343,548,1234,1423,1488,2503,2536,2793,3559,3583,
16,184,340,358,606,647,1402,1618,1727,2807,2895,3090,3863,3887,
120,147,207,231,289,401,1157,1227,2145,2307,2368,2558,3363,3387,
24,70,109,276,990,1043,1745,1786,2123,2767,2775,3203,4259,4283,
4,169,260,456,778,959,1192,2004,2039,2434,2682,3119,4175,4199,
105,177,250,372,435,644,1452,1634,2071,2453,2532,3004,3588,3612,
114,186,259,381,444,629,1461,1643,2080,2462,2541,3013,3597,3621,
42,48,65,190,722,973,1128,1240,2049,2171,2208,2740,3264,3288,
3,66,291,302,329,750,1252,1371,1830,2182,2451,2517,3507,3531,
209,217,283,541,611,1028,1691,1903,1961,2217,2771,2847,3827,3851,
60,169,294,832,838,911,1395,1475,1918,2540,2631,2998,4054,4078,
82,120,156,312,682,880,1605,1916,1960,2816,2982,3040,4096,4120,
5,173,347,353,619,636,1415,1631,1716,2796,2884,3079,3852,3876,
9,130,167,557,573,869,1342,1546,1637,2558,2633,2717,3773,3797,
160,214,228,480,649,837,1139,1729,1752,2346,2809,2851,3865,3889,
85,137,189,193,208,418,1165,1167,1202,2245,2968,3237,3301,3325,
38,61,68,186,742,969,1148,1236,2045,2167,2228,2736,3284,3308,
13,119,191,316,745,1070,1434,1713,1825,2386,2905,3231,3961,3985,
22,143,156,562,570,882,1331,1559,1650,2547,2622,2730,3786,3810,
0,189,256,476,774,955,1188,2000,2035,2430,2678,3115,4171,4195,
79,162,165,216,385,844,1465,2020,2045,2194,2545,2747,3601,3625,
108,180,253,375,438,647,1455,1637,2074,2456,2535,3007,3591,3615,
26,173,289,381,1044,1074,1458,1822,2154,2236,3147,3234,4290,4314,
175,254,345,510,813,912,1544,1992,2112,3015,3072,3143,4128,4152,
90,113,310,322,352,533,1243,1432,1497,2512,2521,2802,3568,3592,
27,99,304,317,471,857,1551,1857,2095,2312,2631,3048,3687,3711,
93,116,289,325,355,536,1246,1435,1500,2515,2524,2805,3571,3595,
57,114,245,271,715,865,1094,1106,1194,2274,2422,2589,3330,3354,
35,46,75,579,588,1013,1308,1532,2093,2248,2824,3173,4229,4253,
93,121,173,192,201,426,1173,1175,1210,2253,2952,3221,3309,3333,
260,342,357,797,896,1019,1248,1561,1877,2297,2957,3138,4013,4037,
124,195,277,316,1005,1057,1742,2007,2085,2291,3165,3179,4221,4245,
26,50,117,281,397,526,1354,1606,1980,2475,2660,2686,3742,3766,
157,159,184,267,354,435,1203,1442,1515,2595,2863,2916,3651,3675,
255,340,353,616,678,1040,1711,1758,1803,2698,2838,3079,3894,3918,
41,64,71,189,721,972,1151,1239,2048,2170,2231,2739,3287,3311,
44,116,297,334,464,850,1544,1850,2088,2305,2624,3065,3680,3704,
127,134,141,220,736,772,1221,1753,1864,2270,2301,3165,3357,3381,
123,150,210,234,292,404,1160,1230,2148,2310,2371,2561,3366,3390,
59,76,77,419,683,945,1499,1671,2119,2448,2579,3097,3635,3659,
250,347,356,811,910,1009,1262,1575,1891,2287,2971,3128,4027,4051,
66,175,300,820,838,893,1401,1481,1900,2522,2637,2980,4036,4060,
88,133,284,339,633,840,1273,1920,2083,2693,2930,3000,4056,4080,
8,129,277,295,451,711,1182,1791,1943,2225,2509,2871,3927,3951,
30,41,94,583,598,1008,1303,1527,2088,2243,2819,3168,4224,4248,
13,59,108,204,223,529,1609,1954,2027,2365,2689,2882,3745,3769,
75,98,295,331,337,542,1228,1417,1506,2497,2530,2787,3553,3577,
22,50,83,167,258,765,1102,1419,1667,2182,2273,3028,3262,4317,
85,123,159,315,685,883,1584,1919,1963,2819,2985,3043,4099,4123,
58,75,76,418,682,944,1498,1670,2118,2471,2578,3096,3634,3658,
169,248,339,504,807,930,1538,2010,2130,3009,3090,3137,4146,4170,
39,61,100,267,1005,1034,1736,1777,2114,2766,2782,3194,4250,4274,
5,126,274,292,448,708,1179,1788,1940,2222,2506,2868,3924,3948,
3,109,181,330,759,1060,1424,1727,1839,2376,2919,3221,3975,3999,
		others => 0);
	end function;

	function init_vector_shifts return vector_shifts is
	begin
		return (
0,3,13,8,11,2,0,0,3,13,0,1,0,0,
1,10,9,0,11,14,0,7,0,4,0,13,0,0,
13,3,5,10,8,0,0,8,13,1,0,4,0,0,
14,0,3,8,12,2,0,0,4,14,0,1,0,0,
12,8,0,10,13,2,1,0,6,12,0,8,0,0,
7,8,8,0,0,5,4,5,0,10,0,8,0,0,
8,4,9,12,8,0,8,11,0,0,4,1,0,0,
14,0,3,8,12,2,0,0,4,14,0,1,0,0,
7,2,10,12,0,2,7,0,8,7,0,14,0,0,
2,14,5,0,8,9,6,0,11,0,14,2,0,0,
0,3,9,8,8,2,13,0,12,0,7,3,0,0,
0,2,8,6,6,10,0,7,12,0,7,3,0,14,
14,4,9,0,2,10,0,10,1,12,0,13,0,0,
2,14,5,0,8,9,6,0,11,0,13,2,0,0,
3,14,2,9,5,0,12,0,7,4,0,4,0,0,
5,9,5,8,12,0,9,11,0,13,2,0,0,0,
10,14,0,3,3,0,9,0,8,3,0,0,0,0,
6,7,8,14,0,4,4,5,0,10,0,8,0,0,
8,0,3,1,12,0,0,7,1,8,0,1,0,0,
1,1,11,11,0,12,14,3,0,5,0,2,0,0,
8,1,1,8,13,0,3,9,0,0,2,0,0,0,
0,0,7,13,2,0,4,7,0,8,11,0,0,0,
3,9,5,12,0,3,0,0,14,0,4,12,0,0,
14,12,0,6,2,11,0,14,8,8,0,9,0,0,
2,0,9,1,7,13,14,3,0,0,14,7,0,0,
6,6,7,5,2,0,2,6,0,0,3,5,0,0,
4,1,13,1,0,1,0,1,8,13,0,6,0,0,
12,2,4,9,8,0,0,7,12,0,0,4,0,0,
12,9,0,13,13,0,13,0,12,3,8,0,0,0,
14,4,9,0,2,10,0,10,1,12,0,13,0,0,
8,0,1,7,13,0,2,8,0,0,1,0,0,0,
10,8,8,7,0,14,1,7,0,11,4,0,0,0,
4,14,0,8,12,2,0,0,4,14,0,1,0,0,
0,11,14,13,1,7,0,4,6,0,1,7,0,0,
3,8,1,13,0,14,11,5,0,3,10,0,0,0,
9,11,7,6,0,10,0,7,7,12,0,9,0,0,
5,2,13,1,0,1,0,1,8,13,0,6,0,0,
7,7,8,0,0,4,4,5,0,10,0,8,0,0,
0,2,9,6,7,11,0,7,13,0,8,3,0,0,
3,12,12,7,10,0,1,2,0,4,0,10,0,0,
5,8,12,12,3,0,0,10,0,9,0,9,0,0,
0,12,0,13,2,7,0,4,6,0,1,7,0,0,
5,2,13,1,0,1,0,1,8,13,0,7,0,0,
11,9,8,7,0,14,1,8,0,12,4,0,0,0,
8,13,3,11,10,0,0,11,0,7,14,0,0,0,
12,8,11,0,13,2,1,0,6,12,0,8,0,0,
2,9,5,11,0,3,0,14,14,0,3,11,0,0,
9,10,4,2,0,2,0,1,12,8,0,3,0,0,
1,3,2,0,7,8,0,1,13,4,0,5,0,0,
8,14,10,12,8,0,8,6,0,13,9,0,0,0,
8,4,9,12,9,0,9,12,0,0,5,1,0,0,
6,7,7,14,0,4,3,4,0,9,0,7,0,0,
2,14,5,0,8,9,6,0,11,0,13,2,0,0,
8,13,3,11,9,0,14,10,0,6,14,0,0,0,
3,14,2,9,5,0,12,0,7,4,0,4,0,0,
9,11,4,2,0,2,0,1,12,8,0,3,0,0,
13,10,0,14,13,0,14,0,12,3,8,0,0,0,
5,2,13,1,0,1,0,1,8,13,0,7,0,0,
5,2,13,1,0,2,0,1,8,13,0,7,0,0,
0,3,9,8,8,2,13,0,11,0,7,3,0,0,
2,14,5,0,8,9,6,0,11,0,13,1,0,0,
13,9,8,5,8,0,7,0,10,1,11,0,0,0,
1,11,9,0,12,0,0,8,1,4,14,0,0,0,
12,7,0,10,12,2,1,0,6,11,0,7,0,0,
9,1,7,9,0,7,11,0,3,7,0,2,0,0,
14,12,0,6,1,11,0,14,8,8,0,9,0,0,
1,11,9,0,12,0,0,8,1,4,14,0,0,0,
10,5,6,9,12,0,10,12,0,13,2,0,0,0,
2,0,7,0,7,3,12,0,9,0,11,13,0,0,
6,5,1,0,13,10,4,14,0,7,0,11,0,0,
4,1,13,0,0,1,0,0,7,12,0,6,0,0,
9,4,0,1,12,1,0,8,2,9,0,1,0,0,
14,12,0,6,2,11,0,14,8,8,0,9,0,0,
13,14,13,8,11,0,4,2,0,7,1,0,0,0,
2,8,0,0,12,14,11,4,0,2,9,0,0,0,
2,8,0,0,12,14,11,4,0,2,9,0,0,0,
0,4,9,8,9,2,13,0,12,0,7,3,0,0,
13,9,8,5,9,0,8,0,11,2,11,0,0,0,
8,7,0,8,0,7,11,0,3,7,0,2,0,0,
2,14,5,0,8,10,6,0,11,0,14,2,0,0,
13,12,9,8,11,0,2,10,0,2,0,9,0,0,
7,7,13,7,0,5,11,0,14,0,11,4,0,0,
14,14,6,12,1,0,3,6,0,7,10,0,0,0,
13,10,0,14,14,0,14,0,13,3,8,0,0,0,
5,5,6,5,1,0,2,6,0,0,2,4,0,0,
8,0,3,1,12,0,0,7,1,8,0,1,0,0,
7,3,9,12,8,0,8,11,0,0,4,1,0,0,
3,12,1,0,2,6,0,7,1,0,3,5,0,0,
12,2,4,9,8,0,0,7,12,0,0,4,0,0,
4,6,0,2,0,12,0,0,13,0,9,7,0,0,
1,0,6,14,6,2,12,0,9,0,10,12,0,0,
8,0,10,12,8,0,8,6,0,13,9,0,0,0,
13,14,13,8,11,0,5,2,0,7,1,0,0,0,
8,0,1,7,13,0,2,8,0,0,2,0,0,0,
8,7,0,8,0,7,11,0,3,7,0,2,0,0,
6,5,1,0,13,9,4,14,0,7,0,11,0,0,
8,13,3,11,9,0,0,10,0,6,14,0,0,0,
8,2,11,12,0,3,8,0,8,8,0,0,0,0,
7,0,0,7,12,0,2,8,0,14,1,0,0,0,
4,8,11,12,3,0,14,9,0,9,0,9,0,0,
5,9,5,9,12,0,9,12,0,13,2,0,0,0,
13,10,0,14,13,0,13,0,12,3,8,0,0,0,
0,2,9,6,7,11,0,7,13,0,8,3,0,0,
13,3,5,10,8,0,0,8,13,1,0,4,0,0,
0,12,0,14,2,8,0,4,7,0,2,8,0,0,
10,5,6,9,12,0,10,12,0,13,2,0,0,0,
9,10,4,2,0,2,0,0,12,8,0,3,0,0,
8,7,0,8,0,7,11,0,3,7,0,2,0,0,
2,14,5,0,8,9,6,0,11,0,13,2,0,0,
9,13,3,11,10,0,0,11,0,7,14,0,0,0,
0,14,7,2,12,0,3,7,0,8,11,0,0,0,
7,0,0,7,12,0,2,8,0,14,1,0,0,0,
12,13,13,8,11,0,4,2,0,7,1,0,0,0,
4,1,13,0,0,1,0,0,7,12,0,6,0,0,
14,10,8,5,9,0,8,0,11,2,11,0,0,0,
3,8,1,13,0,14,12,5,0,3,10,0,0,0,
8,14,10,12,7,0,8,6,0,13,9,0,0,0,
3,8,1,13,0,14,11,5,0,3,10,0,0,0,
0,2,9,6,7,11,0,8,13,0,8,4,0,0,
11,9,8,7,0,14,1,8,0,12,4,0,0,0,
13,3,5,10,9,0,0,8,13,1,0,4,0,0,
6,6,7,5,2,0,2,6,0,0,2,5,0,0,
14,12,0,6,1,11,0,13,8,8,0,9,0,0,
14,10,12,8,11,0,2,10,0,2,0,9,0,0,
2,9,5,12,0,3,0,0,14,0,4,12,0,0,
5,6,1,3,0,13,1,0,14,0,10,8,0,0,
0,2,8,6,7,11,0,7,12,0,8,3,0,0,
3,14,2,9,5,0,12,0,7,4,0,4,0,0,
9,0,3,1,12,0,0,7,1,8,0,1,0,0,
0,3,8,7,8,2,12,0,11,0,6,2,0,0,
8,0,10,12,8,0,8,6,0,14,10,0,0,0,
3,12,2,0,2,7,0,7,1,0,3,5,0,0,
14,12,9,8,11,0,2,10,0,2,0,9,0,0,
8,13,3,11,10,0,0,11,0,7,14,0,0,0,
1,3,2,0,7,8,0,2,13,5,0,6,0,0,
0,12,0,13,2,8,0,4,7,0,1,8,0,0,
4,1,13,0,0,1,0,1,8,13,0,6,0,0,
8,0,1,7,13,0,2,8,0,14,1,0,0,0,
13,9,8,5,9,0,8,0,11,1,11,0,0,0,
2,0,6,14,7,2,12,0,9,0,10,12,0,0,
10,8,8,7,0,14,1,7,0,12,4,0,0,0,
13,9,8,5,9,0,8,0,11,1,11,0,0,0,
2,14,5,0,8,9,6,0,11,0,13,1,0,0,
5,5,6,5,1,0,2,6,0,0,2,4,0,0,
6,6,13,7,0,5,10,0,13,0,11,3,0,0,
14,10,12,9,12,0,2,10,0,3,0,9,0,0,
13,10,0,14,13,0,14,0,12,3,8,0,0,0,
12,8,11,0,13,2,1,0,6,12,0,8,0,0,
14,0,3,8,12,2,0,0,4,14,0,1,0,0,
2,0,6,14,7,2,12,0,9,0,10,12,0,0,
10,11,5,2,0,3,0,1,13,8,0,3,0,0,
3,0,5,0,8,10,6,0,11,0,14,2,0,0,
14,10,9,0,4,8,0,13,3,12,0,3,0,0,
8,11,7,6,0,10,0,7,7,12,0,9,0,0,
9,0,11,12,8,0,8,6,0,14,10,0,0,0,
3,14,2,9,5,0,12,0,7,4,0,4,0,0,
12,2,4,9,8,0,0,7,12,0,0,4,0,0,
8,7,0,8,0,7,11,0,3,7,0,2,0,0,
10,8,8,7,0,14,1,7,0,11,3,0,0,0,
5,5,1,0,13,9,4,14,0,6,0,10,0,0,
0,12,0,13,2,8,0,4,7,0,2,8,0,0,
6,6,13,0,6,4,10,0,13,0,10,3,0,0,
13,9,8,4,8,0,7,0,10,1,10,0,0,0,
12,8,11,0,13,3,2,0,7,12,0,8,0,0,
6,6,7,5,2,0,2,6,0,0,3,5,0,0,
7,7,14,7,0,5,11,0,14,0,11,4,0,0,
5,9,5,8,11,0,9,11,0,13,2,0,0,0,
7,2,10,12,0,3,7,0,8,7,0,0,0,0,
2,1,11,11,0,13,14,4,0,6,0,2,0,0,
13,3,8,0,1,9,0,9,0,11,0,12,0,0,
14,10,12,8,12,0,2,10,0,3,0,9,0,0,
10,5,6,9,12,0,10,12,0,13,2,0,0,0,
6,7,7,14,0,4,3,4,0,9,0,7,0,0,
6,6,13,7,0,4,10,0,13,0,11,3,0,0,
0,12,0,13,2,8,0,4,7,0,1,8,0,0,
14,12,0,6,1,11,0,13,8,8,0,9,0,0,
0,14,7,2,12,0,3,6,0,7,10,0,0,0,
4,14,0,9,12,3,0,1,4,14,0,1,0,0,
9,11,4,2,0,3,0,1,12,8,0,3,0,0,
14,4,9,0,2,9,0,9,1,12,0,13,0,0,
13,0,11,5,1,10,0,13,7,7,0,8,0,0,
2,14,4,0,8,9,5,0,10,0,13,1,0,0,
2,14,5,0,8,9,6,0,10,0,13,1,0,0,
0,10,10,0,4,8,14,0,4,13,0,4,0,0,
8,0,3,1,12,0,0,7,1,8,0,1,0,0,
13,14,13,8,11,0,4,2,0,7,1,0,0,0,
5,9,6,9,12,0,10,12,0,13,2,0,0,0,
8,2,11,12,0,3,8,0,8,8,0,0,0,0,
4,8,11,12,2,0,14,9,0,9,0,8,0,0,
14,10,12,8,12,0,2,10,0,2,0,9,0,0,
10,11,5,3,0,3,0,1,13,8,0,4,0,0,
0,3,9,7,8,2,12,0,11,0,7,2,0,0,
9,11,7,6,0,10,0,7,7,12,0,9,0,0,
4,1,13,0,0,1,0,0,7,12,0,6,0,0,
0,11,14,13,1,7,0,3,6,0,1,7,0,0,
1,0,8,0,7,13,13,3,0,0,14,7,0,0,
4,0,3,10,5,0,13,0,7,5,0,4,0,0,
5,8,12,12,3,0,14,9,0,9,0,9,0,0,
12,7,0,10,12,2,1,0,6,11,0,7,0,0,
3,8,0,13,0,14,11,5,0,3,10,0,0,0,
1,2,1,0,7,8,0,1,13,4,0,5,0,0,
1,10,9,0,11,14,0,7,0,4,0,13,0,0,
0,3,9,7,8,2,12,0,11,0,7,2,0,0,
12,8,0,10,13,2,1,0,6,12,0,8,0,0,
10,13,0,3,2,0,9,0,8,2,0,0,0,0,
8,14,10,12,7,0,8,6,0,13,9,0,0,0,
14,4,9,0,2,9,0,10,1,12,0,13,0,0,
12,7,0,10,12,2,1,0,6,11,0,7,0,0,
8,7,0,8,0,7,11,0,3,7,0,2,0,0,
4,6,0,3,0,13,0,0,14,0,10,7,0,0,
8,0,1,7,13,0,2,8,0,0,2,0,0,0,
10,14,0,3,3,0,9,0,8,2,0,0,0,0,
4,13,13,8,11,0,2,3,0,5,0,11,0,0,
3,12,2,0,2,6,0,7,1,0,3,5,0,0,
3,0,2,9,5,0,12,0,7,5,0,4,0,0,
0,12,0,14,2,8,0,4,7,0,2,8,0,0,
7,8,8,0,0,4,4,5,0,10,0,8,0,0,
4,1,13,0,0,1,0,1,7,12,0,6,0,0,
2,0,7,0,7,3,12,0,9,0,11,13,0,0,
3,12,1,0,2,6,0,7,1,0,3,5,0,0,
6,6,13,7,0,5,10,0,13,0,11,3,0,0,
1,3,2,0,7,8,0,2,13,5,0,6,0,0,
5,5,6,5,1,0,2,6,0,0,2,4,0,0,
4,6,0,2,0,12,0,0,13,0,9,7,0,0,
2,0,6,14,7,3,12,0,9,0,10,12,0,0,
8,1,1,8,13,0,3,9,0,0,2,0,0,0,
4,1,13,0,0,1,0,0,7,12,0,6,0,0,
0,0,7,13,2,0,4,7,0,8,11,0,0,0,
2,9,5,11,0,3,0,0,14,0,4,12,0,0,
3,12,1,0,2,6,0,7,1,0,3,5,0,0,
6,7,8,14,0,4,4,5,0,9,0,7,0,0,
4,6,0,3,0,13,0,0,14,0,10,7,0,0,
0,9,11,2,14,3,0,4,8,0,8,12,0,0,
9,13,3,11,10,0,0,11,0,7,14,0,0,0,
12,7,0,10,12,2,1,0,6,11,0,7,0,0,
9,10,4,2,0,2,0,1,12,8,0,3,0,0,
9,1,7,9,0,8,12,0,3,8,0,3,0,0,
0,14,7,2,12,0,3,7,0,8,11,0,0,0,
2,1,11,11,0,13,14,3,0,5,0,2,0,0,
8,2,11,12,0,3,8,0,8,8,0,0,0,0,
1,10,9,0,12,14,0,7,1,4,0,13,0,0,
9,4,0,1,12,1,0,8,2,9,0,1,0,0,
9,13,14,3,2,0,9,0,7,2,0,0,0,0,
5,5,6,5,2,0,2,6,0,0,2,4,0,0,
6,7,8,14,0,4,4,5,0,10,0,8,0,0,
1,10,9,0,12,0,0,8,1,4,0,13,0,0,
10,11,5,3,0,3,0,1,13,8,0,4,0,0,
10,11,5,2,0,3,0,1,13,8,0,4,0,0,
14,0,3,8,12,2,0,0,4,14,0,1,0,0,
4,14,0,9,12,3,0,0,4,14,0,1,0,0,
14,10,12,8,12,0,2,10,0,2,0,9,0,0,
14,10,9,0,4,8,0,13,3,12,0,3,0,0,
5,2,13,1,0,1,0,1,8,13,0,7,0,0,
13,12,9,8,11,0,2,10,0,2,0,9,0,0,
0,3,9,7,8,2,12,0,11,0,7,3,0,0,
1,3,2,0,7,8,0,1,13,4,0,5,0,0,
8,4,9,12,8,0,8,11,0,0,5,1,0,0,
3,14,2,9,5,0,12,0,7,4,0,4,0,0,
3,12,2,0,2,6,0,7,1,0,3,5,0,0,
2,1,11,12,0,13,14,4,0,6,0,2,0,0,
2,9,5,11,0,3,0,0,14,0,4,11,0,0,
1,11,9,0,12,0,0,8,1,4,14,0,0,0,
5,5,6,5,1,0,2,6,0,0,2,4,0,0,
13,9,8,4,8,0,7,0,10,1,11,0,0,0,
13,9,8,4,8,0,7,0,10,1,11,0,0,0,
2,8,0,13,0,14,11,4,0,3,9,0,0,0,
8,7,10,6,0,10,0,7,7,11,0,8,0,0,
13,10,0,14,13,0,14,0,12,3,8,0,0,0,
6,6,7,5,2,0,2,6,0,0,3,5,0,0,
6,7,7,14,0,4,3,5,0,9,0,7,0,0,
8,2,10,12,0,3,7,0,8,8,0,0,0,0,
2,14,4,0,8,9,5,0,10,0,13,1,0,0,
1,1,11,11,0,12,14,3,0,5,0,1,0,0,
13,9,8,5,9,0,8,0,11,1,11,0,0,0,
10,8,7,0,6,14,0,7,0,11,3,0,0,0,
0,9,11,2,14,3,0,4,8,0,8,12,0,0,
10,9,8,7,0,14,1,8,0,12,4,0,0,0,
10,8,8,0,6,14,0,7,0,11,3,0,0,0,
4,8,11,12,3,0,14,9,0,9,0,9,0,0,
5,5,6,5,1,0,2,6,0,0,2,4,0,0,
13,12,0,6,1,11,0,13,8,8,0,9,0,0,
0,2,8,6,7,11,0,7,12,0,8,3,0,0,
8,14,10,12,7,0,8,6,0,13,9,0,0,0,
8,4,9,12,8,0,9,12,0,0,5,1,0,0,
9,4,5,8,11,0,9,11,0,12,1,0,0,0,
6,7,7,14,0,4,3,4,0,9,0,7,0,0,
0,10,12,3,0,3,5,0,9,0,9,13,0,0,
5,2,13,1,0,1,0,1,8,13,0,7,0,0,
2,0,7,0,7,3,12,0,9,0,11,12,0,0,
6,6,13,7,0,5,10,0,13,0,11,3,0,0,
0,14,7,2,12,0,3,7,0,7,10,0,0,0,
13,9,8,5,9,0,8,0,11,1,11,0,0,0,
12,8,11,0,13,3,1,0,7,12,0,8,0,0,
2,0,8,0,7,13,14,3,0,0,14,7,0,0,
3,0,3,9,5,0,13,0,7,5,0,4,0,0,
8,4,9,12,9,0,9,12,0,0,5,1,0,0,
9,11,7,6,0,11,0,8,8,12,0,9,0,0,
12,8,11,0,13,3,1,0,7,12,0,8,0,0,
8,11,7,6,0,10,0,7,7,12,0,9,0,0,
1,11,9,0,12,0,0,8,1,4,14,0,0,0,
0,2,8,6,6,11,0,7,12,0,7,3,0,0,
3,9,5,12,0,4,0,0,14,0,4,12,0,0,
13,10,0,13,13,0,13,0,12,3,8,0,0,0,
2,0,6,14,7,3,12,0,9,0,11,12,0,0,
3,10,5,12,0,4,0,0,14,0,4,12,0,0,
7,7,13,7,0,5,10,0,13,0,11,3,0,0,
0,9,11,0,2,3,0,4,9,0,8,12,0,0,
6,5,1,0,13,9,4,14,0,6,0,10,0,0,
14,10,12,8,12,0,2,10,0,2,0,9,0,0,
5,1,4,0,13,9,3,13,0,6,0,10,0,0,
14,10,10,0,4,8,0,13,4,13,0,4,0,0,
3,12,2,0,2,6,0,7,1,0,3,5,0,0,
7,7,14,7,0,5,11,0,14,0,11,4,0,0,
4,7,11,12,2,0,14,9,0,9,0,8,0,0,
3,14,2,9,5,0,12,0,7,4,0,4,0,0,
6,7,8,14,0,4,4,5,0,10,0,8,0,0,
8,13,3,11,10,0,0,11,0,7,14,0,0,0,
7,0,0,7,12,0,2,8,0,14,1,0,0,0,
2,9,5,11,0,3,0,0,14,0,4,11,0,0,
0,2,8,6,7,11,0,7,12,0,7,3,0,0,
4,6,0,3,0,12,0,0,13,0,9,7,0,0,
8,11,7,6,0,10,0,7,7,12,0,9,0,0,
0,9,11,2,14,2,0,4,8,0,8,12,0,0,
2,0,7,0,7,3,13,0,10,0,11,13,0,0,
14,10,10,0,4,8,14,0,4,13,0,4,0,0,
0,10,8,0,11,14,0,7,0,4,0,13,0,0,
0,2,8,6,7,11,0,7,12,0,8,3,0,0,
7,2,10,12,0,3,7,0,8,7,0,14,0,0,
13,9,11,8,11,0,2,9,0,2,0,9,0,0,
2,9,5,11,0,3,0,14,14,0,3,11,0,0,
7,0,1,7,12,0,2,8,0,14,1,0,0,0,
13,0,11,5,1,11,0,13,8,8,0,9,0,0,
1,1,11,11,0,12,14,3,0,5,0,1,0,0,
10,8,8,7,0,14,1,7,0,11,4,0,0,0,
6,6,7,5,2,0,2,6,0,0,2,5,0,0,
3,12,12,7,10,0,1,2,0,4,0,10,0,0,
0,3,9,7,7,11,0,8,13,0,8,4,0,0,
2,0,6,14,7,2,12,0,9,0,10,12,0,0,
0,9,12,0,2,3,0,4,9,0,8,13,0,0,
8,1,7,9,0,7,11,0,3,7,0,2,0,0,
3,12,1,0,1,6,0,7,1,0,3,5,0,0,
8,4,13,9,9,0,9,12,0,0,5,1,0,0,
0,2,9,6,7,11,0,7,13,0,8,4,0,0,
7,7,14,7,0,5,11,0,14,0,11,4,0,0,
9,0,10,12,8,0,8,6,0,14,10,0,0,0,
3,8,0,13,0,14,11,5,0,3,10,0,0,0,
8,4,13,9,9,0,9,12,0,0,5,1,0,0,
4,6,0,3,0,12,0,0,14,0,9,7,0,0,
7,0,1,7,12,0,2,8,0,14,1,0,0,0,
1,10,9,0,11,14,0,7,0,4,0,13,0,0,
7,3,9,12,8,0,8,11,0,0,4,0,0,0,
6,6,7,5,2,0,2,6,0,0,2,5,0,0,
9,10,4,2,0,2,0,1,12,8,0,3,0,0,
5,5,7,5,2,0,2,6,0,0,2,4,0,0,
9,13,14,3,2,0,9,0,7,2,0,0,0,0,
5,9,5,9,12,0,9,11,0,13,2,0,0,0,
12,13,13,8,11,0,4,2,0,7,1,0,0,0,
4,0,3,10,5,0,13,0,7,5,0,4,0,0,
13,0,11,5,1,11,0,13,8,8,0,9,0,0,
9,11,7,6,0,10,0,7,8,12,0,9,0,0,
0,3,13,8,11,2,0,0,3,13,0,1,0,0,
2,8,0,0,12,14,11,4,0,3,9,0,0,0,
13,12,9,8,11,0,2,10,0,2,0,9,0,0,
8,11,7,6,0,10,0,7,7,11,0,8,0,0,
1,11,9,0,12,0,0,8,1,4,14,0,0,0,
14,10,9,0,4,8,0,13,3,12,0,3,0,0,
5,8,12,12,3,0,14,9,0,9,0,9,0,0,
0,2,9,6,7,11,0,7,13,0,8,3,0,0,
7,3,12,8,8,0,8,11,0,0,4,0,0,0,
12,13,13,8,10,0,4,2,0,7,1,0,0,0,
8,4,9,12,8,0,8,11,0,0,5,1,0,0,
8,0,3,1,12,0,0,7,1,8,0,1,0,0,
9,4,5,8,11,0,9,11,0,12,1,0,0,0,
13,9,11,8,11,0,2,9,0,2,0,9,0,0,
10,13,0,3,2,0,9,0,8,2,0,0,0,0,
8,7,0,8,0,7,11,0,2,7,0,2,0,0,
3,8,0,13,0,14,11,5,0,3,10,0,0,0,
10,14,0,3,3,0,9,0,8,3,0,0,0,0,
9,10,4,2,0,2,0,1,12,8,0,3,0,0,
13,12,0,5,1,11,0,13,8,8,0,9,0,0,
0,0,7,13,2,0,4,7,0,8,11,0,0,0,
2,1,11,11,0,13,14,4,0,6,0,2,0,0,
2,8,0,0,12,14,11,4,0,3,9,0,0,0,
3,8,0,13,0,14,11,4,0,3,10,0,0,0,
14,4,9,0,1,9,0,9,1,11,0,12,0,0,
12,7,0,10,12,2,1,0,6,12,0,7,0,0,
1,3,2,0,7,8,0,1,13,5,0,6,0,0,
7,7,14,7,0,5,11,0,14,0,11,4,0,0,
3,12,2,0,2,6,0,7,1,0,3,5,0,0,
6,6,13,0,6,4,10,0,13,0,10,3,0,0,
2,8,0,13,0,14,11,4,0,3,10,0,0,0,
13,3,5,10,9,0,0,8,13,1,0,4,0,0,
13,9,8,5,9,0,8,0,11,1,11,0,0,0,
3,12,12,7,10,0,1,2,0,4,0,10,0,0,
1,3,2,0,7,8,0,1,13,5,0,6,0,0,
13,10,0,14,14,0,14,0,13,4,8,0,0,0,
7,8,8,0,0,5,4,5,0,10,0,8,0,0,
3,12,13,8,11,0,1,2,0,5,0,10,0,0,
0,9,11,2,14,3,0,4,8,0,8,12,0,0,
1,1,11,11,0,12,13,3,0,5,0,1,0,0,
1,0,6,14,7,2,12,0,9,0,10,12,0,0,
0,4,9,8,9,2,13,0,12,0,7,3,0,0,
8,0,3,0,12,0,0,7,1,8,0,1,0,0,
4,1,13,0,0,1,0,0,7,12,0,6,0,0,
3,12,1,0,1,6,0,7,1,0,3,5,0,0,
0,3,9,7,8,2,12,0,11,0,7,2,0,0,
2,9,5,11,0,3,0,14,14,0,4,11,0,0,
5,8,12,12,3,0,14,9,0,9,0,9,0,0,
1,1,11,11,0,12,13,3,0,5,0,1,0,0,
14,10,10,0,4,8,0,13,3,13,0,4,0,0,
13,2,5,10,8,0,0,7,12,1,0,4,0,0,
14,10,10,0,4,8,14,0,4,13,0,4,0,0,
8,7,0,8,0,7,11,0,3,7,0,2,0,0,
12,13,13,8,11,0,4,2,0,7,1,0,0,0,
13,14,13,8,11,0,5,2,0,2,7,0,0,0,
3,12,2,0,2,6,0,7,1,0,3,5,0,0,
12,8,11,0,13,2,1,0,6,12,0,8,0,0,
2,8,0,0,12,14,11,4,0,3,9,0,0,0,
5,2,14,1,0,2,0,1,8,13,0,7,0,0,
5,9,5,9,12,0,9,12,0,13,2,0,0,0,
12,2,4,9,8,0,0,7,12,0,0,4,0,0,
0,3,9,7,8,2,12,0,11,0,7,2,0,0,
2,0,7,0,7,3,13,0,10,0,11,13,0,0,
2,12,1,0,1,6,0,7,0,0,3,4,0,0,
8,14,10,12,7,0,8,6,0,13,9,0,0,0,
0,3,13,8,12,2,0,0,4,13,0,1,0,0,
0,3,9,6,7,11,0,8,13,0,8,4,0,0,
13,3,5,10,8,0,0,7,13,1,0,4,0,0,
13,12,0,6,1,11,0,13,8,8,0,9,0,0,
14,10,9,0,4,8,0,13,3,12,0,3,0,0,
8,14,10,12,8,0,8,6,0,13,9,0,0,0,
0,14,7,13,2,0,4,7,0,8,11,0,0,0,
4,6,1,3,0,13,0,0,14,0,10,7,0,0,
14,10,9,0,4,8,0,13,3,12,0,3,0,0,
2,0,9,1,7,13,14,3,0,0,14,7,0,0,
0,9,11,2,14,3,0,4,8,0,8,12,0,0,
9,4,0,1,12,1,0,8,2,9,0,1,0,0,
5,1,4,0,13,9,3,14,0,6,0,10,0,0,
13,12,9,8,11,0,2,10,0,2,0,9,0,0,
8,1,1,8,13,0,2,8,0,0,2,0,0,0,
14,10,9,0,4,8,0,13,3,12,0,3,0,0,
13,14,13,8,11,0,5,2,0,2,7,0,0,0,
14,10,10,0,4,8,14,0,4,13,0,4,0,0,
6,5,1,0,13,9,4,14,0,7,0,11,0,0,
10,8,8,7,0,14,1,7,0,11,3,0,0,0,
13,9,8,5,8,0,7,0,10,1,11,0,0,0,
8,0,6,8,0,7,11,0,2,7,0,2,0,0,
0,9,12,0,2,3,0,4,9,0,8,13,0,0,
5,8,12,12,3,0,14,9,0,9,0,9,0,0,
14,10,9,0,3,8,0,13,3,12,0,3,0,0,
13,3,5,10,8,0,0,8,13,1,0,4,0,0,
3,9,1,13,0,0,12,5,0,3,10,0,0,0,
1,1,11,11,0,12,13,3,0,5,0,1,0,0,
14,4,9,0,1,9,0,9,0,11,0,12,0,0,
6,5,1,0,14,10,4,14,0,7,0,11,0,0,
12,2,4,9,8,0,0,7,12,0,0,4,0,0,
1,3,2,0,7,8,0,1,13,5,0,6,0,0,
0,12,0,13,2,8,0,4,6,0,1,8,0,0,
13,0,11,5,1,11,0,13,8,8,0,9,0,0,
1,0,8,0,7,13,14,3,0,0,14,7,0,0,
3,12,2,0,2,6,0,7,1,0,3,5,0,0,
8,13,3,11,9,0,0,11,0,6,14,0,0,0,
8,14,10,12,8,0,8,6,0,13,9,0,0,0,
2,12,1,0,1,6,0,7,0,0,3,4,0,0,
3,12,12,7,10,0,1,2,0,4,0,10,0,0,
8,13,3,11,9,0,0,10,0,6,14,0,0,0,
3,0,5,0,9,10,6,0,11,0,14,2,0,0,
7,1,10,12,0,2,7,0,8,7,0,14,0,0,
2,14,5,0,8,10,6,0,11,0,14,2,0,0,
1,10,9,0,11,14,0,7,0,4,0,13,0,0,
14,4,9,0,2,10,0,10,1,12,0,13,0,0,
2,9,5,11,0,3,0,14,14,0,4,11,0,0,
0,2,8,6,6,11,0,7,12,0,7,3,0,0,
1,1,11,11,0,12,13,3,0,5,0,1,0,0,
12,2,4,9,8,0,0,7,12,0,0,4,0,0,
13,9,8,5,8,0,7,0,10,1,11,0,0,0,
2,14,5,0,8,10,6,0,11,0,14,2,0,0,
6,5,1,0,13,9,4,14,0,7,0,11,0,0,
13,0,11,5,1,11,0,13,8,8,0,9,0,0,
0,3,8,7,8,1,12,0,11,0,6,2,0,0,
9,13,0,3,2,0,9,0,8,2,0,0,0,0,
6,6,13,7,0,5,10,0,13,0,11,3,0,0,
8,14,10,12,8,0,8,6,0,13,9,0,0,0,
1,3,2,0,7,8,0,1,13,5,0,6,0,0,
14,4,9,0,1,9,0,9,0,11,0,12,0,0,
13,9,7,4,8,0,7,0,10,1,10,0,0,0,
5,8,12,12,3,0,14,9,0,9,0,9,0,0,
6,6,13,7,0,4,10,0,13,0,10,3,0,0,
5,8,12,12,3,0,14,9,0,9,0,9,0,0,
2,8,0,13,0,14,11,4,0,3,10,0,0,0,
9,1,7,9,0,7,11,0,3,8,0,2,0,0,
13,0,11,5,1,10,0,13,7,7,0,8,0,0,
0,12,0,13,2,7,0,4,6,0,1,8,0,0,
1,3,2,0,7,8,0,2,13,5,0,6,0,0,
8,4,9,12,8,0,8,11,0,0,5,1,0,0,
10,8,8,7,0,14,1,7,0,12,4,0,0,0,
0,11,14,13,1,7,0,3,6,0,1,7,0,0,
0,12,0,13,2,8,0,4,7,0,2,8,0,0,
3,8,1,13,0,14,12,5,0,3,10,0,0,0,
0,10,10,0,4,8,14,0,4,13,0,4,0,0,
4,7,11,11,2,0,14,9,0,8,0,8,0,0,
14,4,9,0,2,10,0,10,1,12,0,13,0,0,
13,14,13,8,11,0,4,2,0,7,1,0,0,0,
2,1,11,12,0,13,14,4,0,6,0,2,0,0,
13,9,8,5,9,0,7,0,10,1,11,0,0,0,
0,9,11,0,2,3,0,4,9,0,8,12,0,0,
2,9,5,11,0,3,0,0,14,0,4,11,0,0,
0,3,13,8,11,2,0,0,3,13,0,1,0,0,
1,2,1,0,7,7,0,1,12,4,0,5,0,0,
0,2,8,6,7,11,0,7,12,0,8,3,0,0,
1,11,9,0,12,0,0,8,1,4,14,0,0,0,
3,14,2,9,4,0,12,0,7,4,0,4,0,0,
0,4,9,8,9,2,13,0,12,0,7,3,0,0,
3,12,13,8,11,0,1,2,0,5,0,10,0,0,
2,0,9,1,7,14,14,4,0,0,0,7,0,0,
8,4,13,9,9,0,9,12,0,0,5,1,0,0,
3,0,2,9,5,0,12,0,7,5,0,4,0,0,
1,0,8,0,7,13,14,3,0,0,14,7,0,0,
14,10,10,0,4,8,0,13,3,13,0,4,0,0,
9,4,0,1,12,0,0,8,1,8,0,1,0,0,
3,14,2,9,5,0,12,0,7,5,0,4,0,0,
8,13,3,11,9,0,0,11,0,6,14,0,0,0,
14,10,12,8,11,0,2,10,0,2,0,9,0,0,
8,14,10,12,8,0,8,6,0,13,9,0,0,0,
6,6,13,7,0,4,10,0,13,0,11,3,0,0,
2,1,11,12,0,13,14,4,0,6,0,2,0,0,
4,6,0,3,0,12,0,0,14,0,9,7,0,0,
2,14,5,0,8,9,6,0,11,0,13,2,0,0,
5,9,5,8,12,0,9,11,0,13,2,0,0,0,
2,12,1,0,1,6,0,7,0,0,3,4,0,0,
8,13,3,11,9,0,0,10,0,6,14,0,0,0,
8,4,9,12,8,0,9,12,0,0,5,1,0,0,
0,12,0,13,2,8,0,4,6,0,1,8,0,0,
5,2,13,1,0,1,0,1,8,13,0,7,0,0,
12,2,4,9,8,0,0,7,12,0,0,4,0,0,
14,4,9,0,2,9,0,10,1,12,0,13,0,0,
13,12,0,6,1,11,0,13,8,8,0,9,0,0,
4,1,13,0,0,1,0,1,7,13,0,6,0,0,
14,10,10,0,4,8,0,13,4,13,0,4,0,0,
13,14,13,8,11,0,5,2,0,7,1,0,0,0,
2,12,1,0,1,6,0,7,0,0,3,5,0,0,
5,2,13,1,0,1,0,1,8,13,0,6,0,0,
0,3,13,8,11,2,0,0,3,13,0,1,0,0,
1,3,2,0,7,8,0,1,13,4,0,5,0,0,
0,9,12,0,2,3,0,4,9,0,8,13,0,0,
8,4,9,12,8,0,9,12,0,0,5,1,0,0,
1,11,9,0,12,0,0,8,1,4,14,0,0,0,
0,9,11,2,14,2,0,4,8,0,8,12,0,0,
3,0,5,0,9,10,6,0,11,0,14,2,0,0,
13,9,8,5,9,0,8,0,11,1,11,0,0,0,
10,11,5,2,0,3,0,1,13,8,0,4,0,0,
4,1,13,0,0,1,0,0,7,12,0,6,0,0,
10,14,0,3,2,0,9,0,8,2,0,0,0,0,
14,4,9,0,2,9,0,10,1,12,0,13,0,0,
1,3,2,0,7,8,0,1,13,5,0,6,0,0,
2,9,5,11,0,3,0,14,14,0,4,11,0,0,
6,7,7,14,0,4,3,4,0,9,0,7,0,0,
6,5,1,0,13,9,4,14,0,7,0,11,0,0,
13,9,8,5,9,0,7,0,11,1,11,0,0,0,
2,14,4,0,8,9,5,0,10,0,13,1,0,0,
10,14,0,4,3,0,9,0,8,3,1,0,0,0,
4,6,0,2,0,12,0,0,13,0,9,7,0,0,
2,14,4,0,8,9,5,0,10,0,13,1,0,0,
14,10,12,8,11,0,2,10,0,2,0,9,0,0,
7,7,14,7,0,5,11,0,14,0,11,4,0,0,
2,1,11,11,0,13,14,3,0,5,0,2,0,0,
8,13,2,11,9,0,14,10,0,6,13,0,0,0,
5,7,1,3,0,13,1,0,14,0,10,8,0,0,
2,9,5,11,0,3,0,0,14,0,4,11,0,0,
2,14,5,0,8,10,6,0,11,0,14,2,0,0,
1,2,1,0,7,8,0,1,12,4,0,5,0,0,
14,4,9,0,1,9,0,9,1,12,0,12,0,0,
14,10,8,5,9,0,8,0,11,2,11,0,0,0,
2,9,5,11,0,3,0,14,14,0,3,11,0,0,
4,8,11,12,2,0,14,9,0,9,0,8,0,0,
2,0,8,0,7,13,14,3,0,0,14,7,0,0,
4,7,11,11,2,0,14,9,0,8,0,8,0,0,
8,4,13,9,9,0,9,12,0,0,5,1,0,0,
9,1,7,9,0,7,11,0,3,7,0,2,0,0,
3,8,0,13,0,14,11,5,0,3,10,0,0,0,
6,6,13,0,6,4,10,0,13,0,10,3,0,0,
2,0,6,14,7,2,12,0,9,0,10,12,0,0,
0,2,8,6,6,11,0,7,12,0,7,3,0,0,
0,3,9,8,9,2,13,0,12,0,7,3,0,0,
10,11,5,2,0,3,0,1,13,8,0,3,0,0,
9,14,3,11,10,0,0,11,0,7,14,0,0,0,
13,10,0,14,13,0,14,0,12,3,8,0,0,0,
5,9,5,8,11,0,9,11,0,12,2,0,0,0,
6,7,7,14,0,4,4,5,0,9,0,7,0,0,
14,10,10,0,4,8,14,0,4,13,0,4,0,0,
13,0,11,5,1,11,0,13,7,7,0,9,0,0,
2,14,4,0,8,9,6,0,10,0,13,1,0,0,
0,2,8,6,7,11,0,7,12,0,8,3,0,0,
13,9,8,5,9,0,7,0,11,1,11,0,0,0,
2,0,7,0,7,3,12,0,10,0,11,13,0,0,
14,14,7,2,12,0,3,6,0,7,10,0,0,0,
0,9,12,0,2,3,0,4,9,0,8,13,0,0,
8,2,11,12,0,3,8,0,8,8,0,0,0,0,
9,10,4,2,0,2,0,1,12,8,0,3,0,0,
8,13,2,11,9,0,14,10,0,6,13,0,0,0,
3,12,13,8,11,0,1,2,0,5,0,10,0,0,
5,5,6,5,2,0,2,6,0,0,2,4,0,0,
0,10,10,0,4,8,14,0,4,13,0,4,0,0,
1,1,11,11,0,13,14,3,0,5,0,2,0,0,
9,1,7,9,0,7,11,0,3,8,0,2,0,0,
8,13,3,11,9,0,14,10,0,6,13,0,0,0,
8,13,3,11,9,0,14,10,0,6,14,0,0,0,
4,7,11,11,2,0,14,9,0,8,0,8,0,0,
5,5,6,5,1,0,2,5,0,0,2,4,0,0,
2,9,5,11,0,3,0,14,13,0,3,11,0,0,
14,12,0,6,2,11,0,14,8,8,0,9,0,0,
12,7,0,10,12,2,1,0,6,12,0,8,0,0,
2,0,7,0,7,3,12,0,10,0,11,13,0,0,
2,0,7,0,7,3,12,0,9,0,11,13,0,0,
13,10,0,14,14,0,14,0,13,3,8,0,0,0,
9,1,7,9,0,8,11,0,3,8,0,2,0,0,
13,14,13,8,11,0,4,2,0,7,1,0,0,0,
8,13,2,11,9,0,14,10,0,6,13,0,0,0,
13,3,9,0,1,9,0,9,0,11,0,12,0,0,
3,12,13,8,11,0,1,2,0,5,0,10,0,0,
2,0,5,0,8,10,6,0,11,0,14,2,0,0,
11,9,8,7,0,14,1,8,0,12,4,0,0,0,
12,13,13,8,11,0,4,2,0,7,1,0,0,0,
0,14,7,2,12,0,3,7,0,7,10,0,0,0,
9,4,0,1,12,0,0,7,1,8,0,1,0,0,
4,12,13,8,11,0,2,3,0,5,0,11,0,0,
14,10,10,0,4,8,0,13,3,13,0,4,0,0,
0,11,14,13,1,7,0,4,6,0,1,7,0,0,
6,6,7,5,2,0,2,6,0,0,2,4,0,0,
1,11,9,0,12,0,0,8,1,4,0,13,0,0,
3,12,12,7,10,0,1,2,0,4,0,10,0,0,
14,4,9,0,1,9,0,9,1,11,0,12,0,0,
0,3,13,8,11,2,0,0,3,13,0,1,0,0,
3,0,2,9,5,0,12,0,7,5,0,4,0,0,
4,6,0,3,0,13,0,0,14,0,9,7,0,0,
12,9,14,13,13,0,13,0,12,3,7,0,0,0,
4,14,0,9,12,3,0,0,4,14,0,1,0,0,
13,3,5,10,9,0,0,8,13,1,0,4,0,0,
0,10,10,0,4,8,14,0,4,13,0,4,0,0,
6,7,7,14,0,4,3,4,0,9,0,7,0,0,
12,7,0,10,12,2,1,0,6,12,0,8,0,0,
8,11,7,6,0,10,0,7,7,11,0,8,0,0,
3,0,2,9,5,0,12,0,7,5,0,4,0,0,
0,4,9,8,9,2,13,0,12,0,7,3,0,0,
2,9,5,11,0,3,0,14,13,0,3,11,0,0,
0,12,0,13,2,7,0,4,6,0,1,7,0,0,
10,8,7,0,6,14,0,7,0,11,3,0,0,0,
6,6,13,0,6,4,10,0,13,0,10,3,0,0,
4,6,0,3,0,13,0,0,14,0,9,7,0,0,
1,0,8,0,7,13,13,3,0,0,14,7,0,0,
7,7,13,7,0,5,11,0,14,0,11,4,0,0,
0,3,13,8,12,2,0,0,4,13,0,1,0,0,
9,4,5,8,11,0,9,11,0,12,2,0,0,0,
0,10,12,3,0,3,5,0,9,0,9,13,0,0,
0,4,9,8,9,2,13,0,12,0,7,3,0,0,
2,8,0,13,0,14,11,4,0,3,10,0,0,0,
12,2,4,9,8,0,0,7,12,0,0,4,0,0,
14,14,7,2,12,0,3,6,0,7,10,0,0,0,
9,11,7,6,0,11,0,8,8,12,0,9,0,0,
10,14,0,3,2,0,9,0,8,2,0,0,0,0,
9,1,7,9,0,7,11,0,3,7,0,2,0,0,
7,1,10,11,0,2,7,0,7,7,0,14,0,0,
9,0,11,13,8,0,8,7,0,14,10,0,0,0,
6,5,1,0,13,10,4,14,0,7,0,11,0,0,
5,1,4,0,13,9,3,13,0,6,0,10,0,0,
0,0,7,13,2,0,4,7,0,8,11,0,0,0,
14,10,8,5,9,0,8,0,11,2,11,0,0,0,
9,11,4,2,0,2,0,1,12,8,0,3,0,0,
8,1,1,8,13,0,2,8,0,0,2,0,0,0,
8,10,6,6,0,10,0,7,7,11,0,8,0,0,
1,0,8,0,7,13,13,3,0,0,14,7,0,0,
5,5,6,5,1,0,2,6,0,0,2,4,0,0,
1,0,8,0,7,13,14,3,0,0,14,7,0,0,
8,11,7,6,0,10,0,7,7,11,0,8,0,0,
9,0,11,13,8,0,8,7,0,14,10,0,0,0,
7,3,9,12,8,0,8,11,0,0,4,1,0,0,
4,8,11,12,3,0,14,9,0,9,0,9,0,0,
9,4,0,1,12,0,0,8,1,8,0,1,0,0,
1,3,2,0,7,8,0,1,13,5,0,6,0,0,
10,8,8,7,0,14,1,7,0,11,4,0,0,0,
8,0,6,8,0,7,11,0,2,7,0,2,0,0,
0,11,14,13,1,7,0,3,6,0,1,7,0,0,
0,9,11,2,14,3,0,4,9,0,8,12,0,0,
4,14,0,9,12,3,0,1,4,14,0,1,0,0,
14,4,9,0,1,9,0,9,1,12,0,13,0,0,
0,2,9,6,7,11,0,7,13,0,8,3,0,0,
9,13,0,3,2,0,9,0,8,2,0,0,0,0,
5,9,5,9,12,0,9,11,0,13,2,0,0,0,
0,3,9,7,8,2,13,0,11,0,7,3,0,0,
8,2,10,12,0,3,7,0,8,8,0,0,0,0,
8,11,7,6,0,10,0,7,7,11,0,9,0,0,
1,3,2,0,7,8,0,1,13,5,0,6,0,0,
5,1,4,0,13,9,3,13,0,6,0,10,0,0,
12,9,0,13,13,0,13,0,12,3,8,0,0,0,
13,12,0,6,1,11,0,13,8,8,0,9,0,0,
13,9,8,5,8,0,7,0,10,1,11,0,0,0,
0,0,7,13,2,0,4,7,0,8,11,0,0,0,
8,2,11,12,0,3,8,0,8,8,0,0,0,0,
8,1,1,8,13,0,3,9,0,0,2,0,0,0,
8,7,0,8,0,7,11,0,3,7,0,2,0,0,
0,12,0,13,2,8,0,4,7,0,2,8,0,0,
9,13,0,3,2,0,9,0,7,2,0,0,0,0,
10,8,7,0,6,14,0,7,0,11,3,0,0,0,
14,10,9,0,3,8,0,13,3,12,0,3,0,0,
5,1,4,0,13,9,3,13,0,6,0,10,0,0,
2,0,9,1,7,14,14,4,0,0,0,8,0,0,
0,14,7,2,12,0,3,7,0,7,10,0,0,0,
0,11,14,13,2,7,0,4,6,0,1,7,0,0,
7,3,9,12,8,0,8,11,0,0,4,0,0,0,
14,12,0,6,2,11,0,14,8,8,0,9,0,0,
13,12,9,8,11,0,2,10,0,2,0,9,0,0,
9,10,4,2,0,2,0,1,12,8,0,3,0,0,
3,12,12,8,10,0,1,2,0,4,0,10,0,0,
3,12,13,8,11,0,1,2,0,5,0,10,0,0,
0,10,12,0,2,3,0,4,9,0,8,13,0,0,
1,1,11,11,0,12,13,3,0,5,0,1,0,0,
8,2,11,12,0,3,8,0,8,8,0,0,0,0,
0,10,10,0,4,8,14,0,4,13,0,4,0,0,
4,8,11,12,3,0,14,9,0,9,0,9,0,0,
2,11,1,0,1,6,0,6,0,0,2,4,0,0,
0,4,9,8,9,2,13,0,12,0,7,3,0,0,
8,2,11,12,0,3,8,0,8,8,0,0,0,0,
8,0,1,7,13,0,2,8,0,0,1,0,0,0,
4,6,0,2,0,12,0,0,13,0,9,7,0,0,
9,11,4,2,0,2,0,1,12,8,0,3,0,0,
0,14,7,2,12,0,3,7,0,8,11,0,0,0,
4,7,11,11,2,0,14,9,0,8,0,8,0,0,
13,14,14,9,11,0,5,2,0,2,7,0,0,0,
2,0,7,0,7,3,12,0,9,0,11,13,0,0,
10,14,0,3,3,0,9,0,8,2,0,0,0,0,
13,3,5,10,9,0,0,8,13,1,0,5,0,0,
7,3,9,12,8,0,8,11,0,0,4,0,0,0,
13,10,0,14,13,0,14,0,13,3,8,0,0,0,
12,13,13,8,10,0,4,2,0,1,6,0,0,0,
4,14,0,8,12,2,0,0,4,14,0,1,0,0,
14,0,3,8,12,2,0,0,4,14,0,1,0,0,
0,3,9,8,8,2,13,0,11,0,7,3,0,0,
1,11,9,0,12,0,0,8,1,4,0,13,0,0,
0,3,8,7,8,1,12,0,11,0,6,2,0,0,
4,14,0,9,12,3,0,1,4,14,0,1,0,0,
8,10,6,6,0,10,0,7,7,11,0,8,0,0,
12,9,0,13,13,0,13,0,12,3,8,0,0,0,
12,13,13,8,11,0,4,2,0,7,1,0,0,0,
1,2,2,0,7,8,0,1,13,4,0,5,0,0,
5,8,12,12,3,0,14,10,0,9,0,9,0,0,
8,13,3,11,10,0,0,11,0,7,14,0,0,0,
4,6,0,2,0,12,0,0,13,0,9,7,0,0,
13,10,0,14,13,0,14,0,12,3,8,0,0,0,
10,8,8,7,0,14,1,7,0,12,4,0,0,0,
9,4,0,1,13,1,0,8,2,9,0,2,0,0,
13,12,9,8,11,0,2,10,0,2,0,9,0,0,
10,8,8,7,0,14,1,7,0,11,3,0,0,0,
13,10,0,14,14,0,14,0,13,4,8,0,0,0,
5,8,12,12,3,0,14,9,0,9,0,9,0,0,
8,2,10,12,0,3,7,0,8,8,0,0,0,0,
10,8,8,0,6,14,1,7,0,11,3,0,0,0,
12,8,11,0,13,2,1,0,6,12,0,8,0,0,
2,11,1,0,1,6,0,6,0,0,2,4,0,0,
13,3,8,0,1,9,0,9,0,11,0,12,0,0,
5,5,6,5,1,0,2,6,0,0,2,4,0,0,
9,0,11,12,8,0,8,6,0,14,10,0,0,0,
6,7,8,14,0,4,4,5,0,9,0,7,0,0,
1,10,9,0,12,14,0,7,1,4,0,13,0,0,
2,1,11,11,0,13,14,4,0,6,0,2,0,0,
2,14,4,0,8,9,5,0,10,0,13,1,0,0,
14,12,9,8,11,0,2,10,0,2,0,9,0,0,
12,9,14,13,13,0,13,0,12,3,7,0,0,0,
8,14,10,12,7,0,8,6,0,13,9,0,0,0,
10,14,0,3,2,0,9,0,8,2,0,0,0,0,
7,2,10,12,0,3,7,0,8,7,0,14,0,0,
9,11,5,2,0,3,0,1,12,8,0,3,0,0,
5,8,12,12,3,0,0,10,0,9,0,9,0,0,
14,4,9,0,2,10,0,10,1,12,0,13,0,0,
1,0,10,11,0,12,13,3,0,5,0,1,0,0,
4,7,11,11,2,0,14,9,0,9,0,8,0,0,
2,9,5,11,0,3,0,14,14,0,3,11,0,0,
1,0,8,0,7,13,13,3,0,0,14,7,0,0,
4,0,3,10,5,0,13,0,7,5,0,4,0,0,
8,0,1,7,13,0,2,8,0,0,2,0,0,0,
14,4,9,0,2,10,0,10,1,12,0,13,0,0,
0,9,11,2,14,2,0,4,8,0,8,12,0,0,
9,4,0,1,12,1,0,8,1,9,0,1,0,0,
2,12,1,0,1,6,0,7,0,0,3,5,0,0,
9,1,7,9,0,7,11,0,3,7,0,2,0,0,
8,2,10,12,0,3,7,0,8,8,0,0,0,0,
14,4,9,0,2,10,0,10,1,12,0,13,0,0,
2,9,5,11,0,3,0,14,14,0,3,11,0,0,
0,9,11,2,14,3,0,4,8,0,8,12,0,0,
2,0,9,1,7,14,14,4,0,0,0,8,0,0,
8,2,11,12,0,3,8,0,8,8,0,0,0,0,
8,7,10,6,0,10,0,7,7,11,0,8,0,0,
2,1,11,11,0,13,14,4,0,6,0,2,0,0,
8,11,7,6,0,10,0,7,7,11,0,8,0,0,
5,2,13,1,0,1,0,1,8,13,0,7,0,0,
13,14,14,8,11,0,5,2,0,2,7,0,0,0,
13,9,11,8,11,0,1,9,0,2,0,9,0,0,
8,2,11,12,0,3,8,0,8,8,0,0,0,0,
2,0,9,1,7,14,14,4,0,0,14,7,0,0,
3,0,2,9,5,0,12,0,7,5,0,4,0,0,
12,13,13,8,10,0,4,2,0,1,6,0,0,0,
7,8,8,0,0,5,4,5,0,10,0,8,0,0,
4,14,0,8,12,2,0,0,4,14,0,1,0,0,
5,9,5,8,11,0,9,11,0,12,2,0,0,0,
0,9,11,0,2,3,0,4,9,0,8,12,0,0,
3,9,5,12,0,3,0,0,14,0,4,12,0,0,
7,8,8,0,0,4,4,5,0,10,0,8,0,0,
2,0,9,1,8,14,14,4,0,0,0,8,0,0,
9,4,5,8,11,0,9,11,0,12,1,0,0,0,
10,14,0,4,3,0,9,0,8,3,0,0,0,0,
14,12,0,6,2,11,0,14,8,8,0,9,0,0,
0,2,8,6,7,11,0,7,12,0,8,3,0,0,
2,0,9,1,7,14,14,4,0,0,14,7,0,0,
6,5,1,0,13,9,4,14,0,7,0,11,0,0,
8,11,7,6,0,10,0,7,7,11,0,8,0,0,
8,1,7,8,0,7,11,0,3,7,0,2,0,0,
9,1,7,9,0,7,11,0,3,7,0,2,0,0,
0,9,11,2,14,3,0,4,8,0,8,12,0,0,
2,0,7,0,7,3,12,0,10,0,11,13,0,0,
1,0,8,0,7,13,14,3,0,0,14,7,0,0,
8,0,1,7,13,0,2,8,0,0,2,0,0,0,
8,14,10,12,8,0,8,6,0,13,9,0,0,0,
11,9,8,7,0,14,1,8,0,12,4,0,0,0,
3,8,1,13,0,14,11,5,0,3,10,0,0,0,
13,13,13,8,11,0,4,2,0,7,1,0,0,0,
6,6,7,5,2,0,2,6,0,0,2,5,0,0,
4,1,13,1,0,1,0,1,8,13,0,6,0,0,
9,10,4,2,0,2,0,0,12,8,0,3,0,0,
10,14,0,4,3,0,10,0,8,3,1,0,0,0,
12,8,11,0,13,2,1,0,6,12,0,8,0,0,
6,7,8,14,0,4,4,5,0,10,0,8,0,0,
9,4,5,8,11,0,9,11,0,12,1,0,0,0,
9,10,4,2,0,2,0,0,12,7,0,3,0,0,
8,0,1,7,13,0,2,8,0,0,2,0,0,0,
7,2,10,12,0,3,7,0,8,8,0,0,0,0,
0,3,8,7,8,1,12,0,11,0,6,2,0,0,
3,12,12,7,10,0,1,2,0,4,0,10,0,0,
0,9,11,2,14,3,0,4,8,0,8,12,0,0,
12,8,11,0,13,2,1,0,6,12,0,8,0,0,
3,12,2,0,2,7,0,7,1,0,3,5,0,0,
3,9,1,13,0,14,12,5,0,3,10,0,0,0,
1,11,9,0,12,0,0,8,1,4,0,13,0,0,
8,2,11,12,0,3,7,0,8,8,0,0,0,0,
1,10,9,0,11,14,0,7,1,4,0,13,0,0,
8,13,3,11,9,0,0,10,0,6,14,0,0,0,
12,13,13,8,10,0,4,1,0,1,6,0,0,0,
10,13,0,3,2,0,9,0,8,2,0,0,0,0,
13,2,4,9,8,0,0,7,12,1,0,4,0,0,
1,2,1,0,7,8,0,1,12,4,0,5,0,0,
8,11,7,6,0,10,0,7,7,11,0,8,0,0,
8,14,10,12,7,0,8,6,0,13,9,0,0,0,
2,0,5,0,8,10,6,0,11,0,14,2,0,0,
13,3,5,10,9,0,0,8,13,1,0,4,0,0,
13,14,13,8,11,0,4,2,0,7,1,0,0,0,
8,10,6,5,0,10,0,7,7,11,0,8,0,0,
0,11,14,13,1,7,0,3,6,0,1,7,0,0,
12,2,4,9,8,0,0,7,12,0,0,4,0,0,
12,9,0,13,13,0,13,0,12,3,8,0,0,0,
9,0,11,12,8,0,8,7,0,14,10,0,0,0,
9,4,0,1,12,1,0,8,1,8,0,1,0,0,
8,13,3,11,10,0,0,11,0,7,14,0,0,0,
10,14,0,3,3,0,9,0,8,2,0,0,0,0,
13,9,8,5,9,0,8,0,11,1,11,0,0,0,
0,0,7,13,2,0,4,7,0,8,11,0,0,0,
12,10,0,13,13,0,13,0,12,3,8,0,0,0,
0,2,9,6,7,11,0,7,13,0,8,3,0,0,
8,7,0,8,0,7,11,0,3,7,0,2,0,0,
6,7,7,14,0,4,3,4,0,9,0,7,0,0,
10,8,8,7,0,14,1,7,0,11,3,0,0,0,
9,4,0,1,12,1,0,8,2,9,0,1,0,0,
6,6,7,5,2,0,2,6,0,0,2,5,0,0,
9,4,0,1,12,1,0,8,1,9,0,1,0,0,
4,12,13,8,11,0,2,2,0,5,0,11,0,0,
5,9,6,9,12,0,10,12,0,13,2,0,0,0,
0,14,7,2,12,0,3,7,0,7,10,0,0,0,
4,0,3,10,5,0,13,0,7,5,0,4,0,0,
8,11,7,6,0,10,0,7,7,11,0,8,0,0,
7,2,10,12,0,3,7,0,8,8,0,0,0,0,
1,2,1,0,7,7,0,1,12,4,0,5,0,0,
5,2,13,1,0,1,0,1,8,13,0,6,0,0,
3,10,5,12,0,4,0,0,14,0,4,12,0,0,
5,8,12,12,3,0,14,10,0,9,0,9,0,0,
8,13,3,11,9,0,14,10,0,6,13,0,0,0,
2,0,8,1,7,13,14,3,0,0,14,7,0,0,
0,12,0,13,2,8,0,4,6,0,1,8,0,0,
10,14,0,3,3,0,9,0,8,2,0,0,0,0,
9,4,5,8,11,0,9,11,0,12,1,0,0,0,
12,8,11,0,13,2,1,0,6,12,0,8,0,0,
14,10,12,9,12,0,2,10,0,3,0,10,0,0,
9,4,0,1,12,0,0,8,1,8,0,1,0,0,
14,4,9,0,2,9,0,10,1,12,0,13,0,0,
3,12,13,8,11,0,1,2,0,5,0,11,0,0,
4,12,13,8,11,0,2,2,0,5,0,11,0,0,
9,11,4,2,0,2,0,1,12,8,0,3,0,0,
13,10,0,14,13,0,14,0,13,3,8,0,0,0,
9,4,0,1,12,1,0,8,2,9,0,2,0,0,
4,6,0,3,0,12,0,0,14,0,9,7,0,0,
0,10,8,0,11,14,0,7,0,4,0,13,0,0,
9,11,7,6,0,11,0,8,8,12,0,9,0,0,
1,0,6,14,6,2,12,0,9,0,10,12,0,0,
14,10,10,0,4,8,0,13,3,12,0,4,0,0,
0,14,7,2,12,0,3,7,0,8,11,0,0,0,
14,14,7,2,12,0,3,6,0,7,10,0,0,0,
3,0,3,9,5,0,12,0,7,5,0,4,0,0,
6,5,1,0,14,10,4,14,0,7,0,11,0,0,
14,10,12,9,12,0,2,10,0,3,0,9,0,0,
6,7,8,14,0,4,4,5,0,10,0,8,0,0,
8,14,10,12,8,0,8,6,0,13,9,0,0,0,
0,10,8,0,11,14,0,7,0,3,0,13,0,0,
12,13,13,8,11,0,4,2,0,7,1,0,0,0,
1,1,11,11,0,12,14,3,0,5,0,1,0,0,
12,2,4,9,8,0,0,7,12,0,0,4,0,0,
2,9,5,11,0,3,0,14,14,0,4,11,0,0,
0,4,9,8,9,2,13,0,12,0,7,3,0,0,
2,1,11,11,0,13,14,4,0,6,0,2,0,0,
4,6,0,3,0,13,0,0,14,0,9,7,0,0,
2,0,9,1,7,13,14,3,0,0,14,7,0,0,
8,4,9,12,8,0,8,11,0,0,5,1,0,0,
4,14,0,9,12,3,0,0,4,14,0,1,0,0,
1,11,9,0,12,0,0,8,1,4,14,0,0,0,
12,8,0,10,13,2,1,0,6,12,0,8,0,0,
9,10,4,2,0,2,0,0,12,7,0,3,0,0,
14,12,0,6,2,11,0,14,8,8,0,9,0,0,
8,0,10,12,8,0,8,6,0,14,9,0,0,0,
4,6,1,3,0,13,0,0,14,0,10,7,0,0,
0,3,9,6,7,11,0,8,13,0,8,4,0,0,
9,4,5,8,11,0,9,11,0,12,1,0,0,0,
3,12,12,8,10,0,1,2,0,4,0,10,0,0,
12,2,4,9,8,0,0,7,12,0,0,4,0,0,
14,10,12,8,12,0,2,10,0,2,0,9,0,0,
8,7,10,6,0,10,0,7,7,11,0,8,0,0,
7,0,0,7,12,0,2,8,0,14,1,0,0,0,
9,13,0,3,2,0,9,0,8,2,0,0,0,0,
0,12,0,13,2,7,0,4,6,0,1,7,0,0,
0,10,9,0,11,14,0,7,0,4,0,13,0,0,
1,3,2,0,7,8,0,2,13,5,0,6,0,0,
0,3,8,7,8,2,12,0,11,0,6,2,0,0,
5,1,4,0,13,9,4,14,0,6,0,10,0,0,
6,5,7,5,2,0,2,6,0,0,2,4,0,0,
0,3,9,7,8,2,12,0,11,0,7,2,0,0,
6,7,8,14,0,4,4,5,0,10,0,8,0,0,
6,6,7,5,2,0,2,6,0,0,3,5,0,0,
6,5,1,0,13,9,4,14,0,7,0,11,0,0,
6,7,13,7,0,5,10,0,13,0,11,3,0,0,
1,0,8,0,7,13,14,3,0,0,14,7,0,0,
9,4,0,1,12,1,0,8,1,8,0,1,0,0,
2,0,7,0,7,3,12,0,10,0,11,13,0,0,
4,6,1,3,0,13,1,0,14,0,10,7,0,0,
0,12,0,13,2,8,0,4,6,0,1,8,0,0,
2,12,1,0,1,6,0,7,0,0,3,4,0,0,
14,0,3,8,12,2,0,0,4,14,0,1,0,0,
6,6,13,0,6,4,10,0,13,0,10,3,0,0,
13,9,8,4,8,0,7,0,10,1,11,0,0,0,
2,9,5,11,0,3,0,14,14,0,4,11,0,0,
3,8,0,13,0,14,11,5,0,3,10,0,0,0,
1,3,2,0,7,8,0,1,13,5,0,6,0,0,
3,12,12,8,10,0,1,2,0,4,0,10,0,0,
4,0,3,10,5,0,13,0,7,5,0,4,0,0,
2,0,6,14,7,2,12,0,9,0,10,12,0,0,
8,0,1,7,13,0,2,8,0,0,2,0,0,0,
7,3,9,12,8,0,8,11,0,0,4,0,0,0,
0,3,8,7,8,2,12,0,11,0,6,2,0,0,
2,1,11,11,0,13,14,3,0,5,0,2,0,0,
3,12,1,0,2,6,0,7,1,0,3,5,0,0,
0,10,10,0,4,8,14,0,4,13,0,4,0,0,
6,5,7,5,2,0,2,6,0,0,2,4,0,0,
8,13,3,11,10,0,0,11,0,7,14,0,0,0,
4,0,3,9,5,0,13,0,7,5,0,4,0,0,
4,8,12,12,3,0,14,9,0,9,0,9,0,0,
12,8,11,0,13,2,1,0,6,12,0,8,0,0,
2,14,5,0,8,9,6,0,11,0,13,2,0,0,
0,14,7,2,12,0,3,6,0,7,10,0,0,0,
14,12,0,6,2,11,0,14,8,8,0,9,0,0,
9,0,11,13,8,0,8,7,0,14,10,0,0,0,
7,7,14,7,0,5,11,0,14,0,11,4,0,0,
8,4,9,12,8,0,9,12,0,0,5,1,0,0,
8,1,1,8,13,0,3,9,0,0,2,0,0,0,
3,12,1,0,2,6,0,7,1,0,3,5,0,0,
9,13,14,3,2,0,9,0,7,2,0,0,0,0,
6,5,1,0,13,9,4,14,0,6,0,11,0,0,
5,9,5,8,11,0,9,11,0,13,2,0,0,0,
1,2,1,0,7,8,0,1,13,4,0,5,0,0,
8,2,11,12,0,3,8,0,8,8,0,0,0,0,
6,7,8,14,0,4,4,5,0,10,0,8,0,0,
6,2,5,0,14,10,4,14,0,7,0,11,0,0,
2,0,7,0,7,3,12,0,9,0,11,13,0,0,
9,4,0,1,12,1,0,8,2,9,0,1,0,0,
10,14,0,3,2,0,9,0,8,2,0,0,0,0,
2,11,1,0,1,6,0,7,0,0,2,4,0,0,
14,12,0,6,2,11,0,14,8,8,0,9,0,0,
14,14,7,2,12,0,3,6,0,7,10,0,0,0,
3,12,13,8,11,0,1,2,0,5,0,10,0,0,
0,2,9,6,7,11,0,7,13,0,8,3,0,0,
12,7,0,10,12,2,1,0,6,12,0,8,0,0,
2,9,5,11,0,3,0,0,14,0,4,11,0,0,
2,0,9,1,7,13,14,4,0,0,14,7,0,0,
3,12,13,8,11,0,1,2,0,5,0,10,0,0,
4,6,0,3,0,13,0,0,14,0,9,7,0,0,
8,0,1,7,13,0,2,8,0,14,1,0,0,0,
3,12,12,7,10,0,1,2,0,4,0,10,0,0,
3,14,2,9,4,0,12,0,7,4,0,4,0,0,
2,0,8,1,7,13,14,3,0,0,14,7,0,0,
0,11,14,13,2,7,0,4,6,0,1,7,0,0,
8,7,0,8,0,7,11,0,3,7,0,2,0,0,
9,11,5,2,0,3,0,1,12,8,0,3,0,0,
14,0,3,8,12,2,0,0,4,14,0,1,0,0,
0,9,11,2,14,3,0,4,8,0,8,12,0,0,
1,11,9,0,12,0,0,8,1,4,0,13,0,0,
0,11,14,13,2,7,0,4,6,0,1,7,0,0,
14,10,12,8,12,0,2,10,0,3,0,9,0,0,
13,10,0,14,13,0,14,0,13,3,8,0,0,0,
13,3,5,10,9,0,0,8,13,1,0,4,0,0,
7,7,13,7,0,5,10,0,14,0,11,3,0,0,
6,5,1,0,13,9,4,14,0,6,0,10,0,0,
5,1,4,0,13,9,4,14,0,6,0,10,0,0,
5,9,5,9,12,0,9,12,0,13,2,0,0,0,
13,10,0,14,13,0,14,0,13,3,8,0,0,0,
13,12,9,8,11,0,2,10,0,2,0,9,0,0,
14,12,0,6,1,11,0,13,8,8,0,9,0,0,
10,8,7,0,6,14,0,7,0,11,3,0,0,0,
0,2,9,6,7,11,0,7,13,0,8,3,0,0,
10,8,7,0,6,14,0,7,0,11,3,0,0,0,
6,6,13,0,6,4,10,0,13,0,10,3,0,0,
9,4,5,8,11,0,9,11,0,12,1,0,0,0,
4,12,13,8,11,0,2,2,0,5,0,11,0,0,
3,12,12,7,10,0,1,2,0,4,0,10,0,0,
12,8,0,10,12,2,1,0,6,12,0,8,0,0,
4,6,0,3,0,12,0,0,14,0,9,7,0,0,
8,4,13,9,9,0,9,12,0,0,5,1,0,0,
2,0,6,14,7,2,12,0,9,0,10,12,0,0,
13,13,13,8,11,0,4,2,0,7,1,0,0,0,
9,14,3,12,10,0,0,11,0,7,14,0,0,0,
14,4,9,0,2,9,0,10,1,12,0,13,0,0,
14,4,9,0,2,10,0,10,1,12,0,13,0,0,
8,0,3,0,12,0,0,7,1,8,0,1,0,0,
12,7,0,10,12,2,1,0,6,11,0,7,0,0,
9,11,4,2,0,2,0,1,12,8,0,3,0,0,
3,9,1,13,0,14,12,5,0,3,10,0,0,0,
8,1,1,8,13,0,2,8,0,0,2,0,0,0,
8,4,9,12,8,0,8,11,0,0,5,1,0,0,
10,8,7,0,6,14,0,7,0,11,3,0,0,0,
7,1,10,12,0,2,7,0,8,7,0,14,0,0,
0,9,11,0,2,3,0,4,9,0,8,12,0,0,
9,4,0,1,12,1,0,8,2,9,0,2,0,0,
1,0,10,11,0,12,13,3,0,5,0,1,0,0,
10,8,8,7,0,14,1,7,0,12,4,0,0,0,
9,13,3,11,10,0,0,11,0,7,14,0,0,0,
8,10,6,6,0,10,0,7,7,11,0,8,0,0,
14,4,9,0,2,9,0,10,1,12,0,13,0,0,
9,0,11,12,8,0,8,6,0,14,10,0,0,0,
3,14,2,9,4,0,12,0,7,4,0,3,0,0,
4,6,0,3,0,13,0,0,14,0,10,7,0,0,
5,2,13,1,0,1,0,1,8,13,0,7,0,0,
4,6,1,3,0,13,0,0,14,0,10,7,0,0,
2,0,9,1,7,14,14,4,0,0,14,7,0,0,
14,14,7,2,12,0,3,6,0,7,10,0,0,0,
0,10,12,3,0,3,0,4,9,0,9,13,0,0,
5,1,4,0,13,9,4,14,0,6,0,10,0,0,
7,8,8,0,0,5,4,5,0,10,0,8,0,0,
14,10,8,5,9,0,8,0,11,2,11,0,0,0,
5,5,6,5,1,0,2,6,0,0,2,4,0,0,
8,7,0,8,0,7,11,0,3,7,0,2,0,0,
9,4,0,1,13,1,0,8,2,9,0,2,0,0,
4,1,13,0,0,1,0,1,8,13,0,6,0,0,
4,14,0,9,12,3,0,1,4,14,0,1,0,0,
2,0,6,14,7,2,12,0,9,0,10,12,0,0,
1,3,2,0,7,8,0,1,13,5,0,6,0,0,
6,5,1,0,13,10,4,14,0,7,0,11,0,0,
2,8,0,0,12,14,11,4,0,3,9,0,0,0,
9,13,14,3,2,0,9,0,7,2,0,0,0,0,
13,10,0,14,13,0,14,0,12,3,8,0,0,0,
14,14,6,12,1,0,3,6,0,7,10,0,0,0,
12,2,4,9,8,0,0,7,12,0,0,4,0,0,
4,6,0,2,0,12,0,0,13,0,9,7,0,0,
0,3,9,6,7,11,0,8,13,0,8,4,0,0,
8,1,1,8,13,0,3,8,0,0,2,0,0,0,
1,3,2,0,7,8,0,1,13,4,0,6,0,0,
4,0,3,10,5,0,13,0,7,5,0,4,0,0,
12,13,13,8,10,0,4,2,0,1,6,0,0,0,
13,10,0,14,13,0,14,0,12,3,8,0,0,0,
2,1,11,11,0,13,14,3,0,6,0,2,0,0,
		others => 0);
	end function;
end package body;
