-- code table generated from table_vector.txt by generate_table_vector_vhd.cc
--
-- Copyright 2019 Ahmet Inan <inan@aicodix.de>

use work.ldpc_scalar.all;
use work.ldpc_vector.all;

package table_vector is
	function init_vector_parities return vector_parities;
	function init_vector_counts return vector_counts;
	function init_vector_offsets return vector_offsets;
	function init_vector_shifts return vector_shifts;
end package;

package body table_vector is
	function init_vector_parities return vector_parities is
	begin
		return 270;
	end function;

	function init_vector_counts return vector_counts is
	begin
		return (
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
		others => count_scalar'low);
	end function;

	function init_vector_offsets return vector_offsets is
	begin
		return (
4,5,66,77,79,241,366,405,511,621,726,781,1045,1051,
21,31,47,48,51,102,291,293,304,561,738,809,825,831,
1,2,69,74,82,244,369,402,514,618,729,784,1048,1054,
4,46,88,88,150,161,352,406,431,701,723,768,965,971,
11,44,76,90,261,267,363,451,537,559,786,807,1071,1077,
21,30,67,86,158,215,318,485,516,676,733,755,1019,1025,
6,45,77,91,262,268,364,452,538,560,787,808,1072,1078,
18,34,44,48,51,105,288,290,301,558,741,806,822,828,
33,50,66,81,248,264,433,500,518,574,788,796,1052,1058,
5,30,70,76,112,174,297,444,482,554,628,714,978,984,
6,12,25,69,101,128,338,398,496,619,660,668,932,938,
1,16,72,73,81,190,314,343,460,542,613,625,877,883,
7,29,56,65,74,78,335,378,471,598,601,605,869,875,
10,43,75,95,260,266,362,450,536,558,791,806,1070,1076,
11,14,24,36,54,177,324,342,526,594,653,667,858,864,
26,49,50,60,76,126,320,335,539,581,590,696,854,860,
22,27,74,80,86,135,311,356,373,626,635,700,890,896,
19,24,77,83,89,132,308,359,376,629,632,697,893,899,
1,17,20,38,63,186,271,354,416,541,566,757,811,1074,
31,51,64,124,162,229,281,394,447,664,680,793,928,934,
5,30,37,139,143,217,330,384,409,640,655,679,943,949,
4,35,69,75,111,179,296,449,481,553,627,719,983,989,
43,62,87,126,201,228,386,498,528,753,768,785,1032,1038,
10,13,29,41,59,176,329,347,525,599,652,666,863,869,
27,64,71,83,83,248,319,353,410,623,646,661,887,893,
8,47,73,93,258,264,360,454,534,562,789,804,1068,1074,
10,15,16,44,180,245,286,308,511,543,556,686,820,826,
53,55,67,133,155,254,425,475,491,555,695,711,959,965,
51,59,71,137,153,252,423,479,489,553,693,709,957,963,
23,28,75,81,87,136,306,357,374,627,630,701,891,897,
1,32,66,72,108,176,299,446,484,556,624,716,980,986,
10,19,43,54,238,243,280,372,497,550,681,778,814,820,
26,44,63,95,110,157,365,409,516,616,635,753,899,905,
3,57,68,144,163,230,414,472,483,684,747,803,948,954,
2,24,42,83,188,267,355,430,458,599,728,808,992,998,
33,36,48,54,76,98,290,306,534,576,589,641,840,846,
11,29,72,79,119,211,389,467,525,580,659,764,923,929,
24,42,61,93,108,161,363,413,520,614,633,751,897,903,
37,39,46,69,84,111,303,362,381,651,715,726,915,921,
3,12,74,75,83,186,316,345,456,544,615,627,879,885,
26,63,70,82,82,247,318,352,409,622,645,660,886,892,
19,38,41,62,122,185,394,422,455,550,725,756,989,995,
44,57,80,85,118,203,284,314,401,584,650,741,848,854,
7,14,20,51,102,194,274,420,464,718,734,762,998,1004,
0,16,29,53,54,132,402,489,508,588,672,721,936,942,
11,15,24,71,251,262,436,447,532,690,692,802,1066,1072,
8,58,76,79,88,225,326,461,495,610,765,801,1029,1035,
1,46,65,117,193,236,295,501,506,607,669,776,1040,1046,
36,38,45,68,89,110,302,361,380,650,714,731,914,920,
4,43,62,114,196,239,298,498,509,610,666,779,1043,1049,
21,37,40,64,124,181,390,424,451,546,721,758,985,991,
6,56,74,83,86,223,324,459,493,608,763,799,1027,1033,
10,14,29,70,250,261,435,446,531,691,695,801,1065,1071,
8,24,57,60,75,79,330,379,472,599,600,602,864,870,
61,86,87,152,172,258,431,442,451,674,712,773,976,982,
39,51,59,125,162,206,286,432,443,587,702,708,966,972,
0,54,71,147,166,233,417,469,480,687,744,800,951,957,
20,25,72,78,84,133,309,354,377,624,633,698,888,894,
2,47,60,118,194,237,296,502,507,608,670,777,1041,1047,
22,31,68,87,159,210,319,480,517,677,734,750,1014,1020,
50,58,70,136,152,257,422,478,488,552,692,708,956,962,
20,35,66,85,157,214,323,484,521,675,732,754,1018,1024,
9,27,76,83,117,215,387,465,523,578,657,762,921,927,
37,41,44,67,88,109,301,360,379,649,719,730,913,919,
6,24,73,80,114,212,384,462,526,581,654,765,918,924,
0,30,52,66,94,138,336,340,342,585,606,736,870,876,
3,25,43,78,189,268,356,431,459,594,729,809,993,999,
22,38,41,65,125,182,391,425,452,547,722,759,986,992,
33,53,60,120,164,231,277,390,449,660,682,795,924,930,
36,48,56,122,165,209,283,435,440,584,705,711,969,975,
28,65,66,78,78,249,320,348,411,618,647,662,882,888,
9,16,22,53,104,196,270,422,466,714,736,764,1000,1006,
42,61,86,131,200,233,385,503,533,752,773,784,1037,1043,
18,32,38,80,168,216,401,478,486,706,746,756,1020,1026,
1,31,53,67,95,139,337,341,343,586,607,737,871,877,
63,85,88,198,225,252,313,392,468,570,738,781,1002,1008,
22,36,39,57,100,211,370,505,512,547,640,686,904,910,
14,19,20,104,170,234,374,414,532,615,644,778,908,914,
1,17,24,48,55,133,403,490,509,589,673,722,937,943,
45,58,81,86,119,198,285,315,396,585,651,742,849,855,
32,33,34,59,185,197,304,440,467,567,574,790,838,844,
17,26,61,69,177,219,274,280,296,566,600,647,830,836,
6,16,25,66,246,263,437,448,533,691,693,803,1067,1073,
9,14,15,43,185,244,285,307,510,542,555,685,819,825,
3,33,49,69,91,141,337,339,345,582,609,733,873,879,
46,59,82,87,114,199,286,316,397,586,652,743,850,856,
16,21,22,106,172,236,376,416,528,617,646,774,910,916,
4,13,75,76,78,187,317,346,457,545,616,628,880,886,
10,17,23,48,105,197,271,423,467,715,737,765,1001,1007,
9,18,42,59,237,242,279,377,496,549,680,777,813,819,
46,65,84,129,198,231,389,501,531,750,771,782,1035,1041,
0,31,71,77,113,175,298,445,483,555,629,715,979,985,
23,37,40,58,101,212,371,506,513,548,641,687,905,911,
22,32,42,49,52,103,288,292,305,562,739,804,826,832,
15,20,21,105,171,235,375,415,533,616,645,779,909,915,
8,14,27,71,97,130,340,400,492,621,662,670,934,940,
34,48,61,121,165,232,278,391,444,661,683,796,925,931,
0,16,19,37,62,191,270,359,415,540,565,756,810,1079,
3,13,22,40,65,188,273,356,418,543,568,759,813,1076,
5,59,70,146,165,232,416,468,485,686,749,799,950,956,
61,86,89,202,223,256,317,390,472,574,742,785,1006,1012,
48,56,68,134,150,255,420,476,486,556,690,712,954,960,
13,28,63,71,179,221,270,276,298,568,602,643,832,838,
18,38,41,59,96,213,366,507,514,549,636,688,900,906,
62,87,88,153,173,259,426,443,452,675,713,768,977,983,
52,54,66,132,154,253,424,474,490,554,694,710,958,964,
11,17,24,68,100,127,337,397,495,618,665,667,931,937,
7,8,18,144,147,254,327,383,524,559,703,794,1058,1064,
41,53,55,121,164,208,282,434,439,583,704,710,968,974,
5,35,51,71,93,143,339,341,347,584,611,735,875,881,
30,31,32,57,183,195,302,438,465,565,572,788,836,842,
12,43,72,208,208,227,351,371,478,632,657,748,1012,1018,
7,17,26,67,247,258,432,449,528,692,694,798,1062,1068,
9,42,74,94,259,265,361,455,535,563,790,805,1069,1075,
40,52,54,120,163,207,287,433,438,582,703,709,967,973,
5,14,76,77,79,188,312,347,458,540,617,629,881,887,
12,18,23,102,168,238,372,418,530,613,642,776,906,912,
4,34,50,70,92,142,338,340,346,583,610,734,874,880,
1,32,39,139,141,219,332,386,411,636,657,681,945,951,
6,15,25,37,55,178,325,343,527,595,648,668,859,865,
64,84,89,155,169,261,428,439,454,677,709,770,973,979,
60,85,86,151,171,263,430,441,450,673,711,772,975,981,
47,54,83,88,115,200,287,317,398,587,653,738,851,857,
17,42,77,207,207,226,350,370,477,631,656,747,1011,1017,
30,39,51,57,73,101,293,309,537,579,592,638,843,849,
5,15,28,52,59,137,407,488,507,593,677,720,941,947,
8,26,75,82,116,214,386,464,522,577,656,767,920,926,
21,35,41,83,171,219,398,475,489,703,749,759,1023,1029,
7,25,74,81,115,213,385,463,527,576,655,766,919,925,
11,16,17,45,181,240,287,309,512,544,557,687,821,827,
32,52,65,125,163,230,276,395,448,665,681,794,929,935,
62,84,87,203,224,257,312,391,473,575,743,780,1007,1013,
11,12,18,49,106,192,272,424,462,716,732,766,996,1002,
22,30,36,78,172,220,399,476,490,704,744,760,1024,1030,
35,52,68,83,250,266,435,502,520,570,790,792,1054,1060,
2,12,25,49,56,134,404,491,504,590,674,723,938,944,
19,36,39,54,97,214,367,508,515,550,637,689,901,907,
17,22,23,107,173,237,377,417,529,612,647,775,911,917,
31,40,52,58,74,96,288,310,538,580,593,639,844,850,
2,32,48,68,90,140,336,338,344,587,608,732,872,878,
1,29,47,82,187,266,354,429,457,598,727,807,991,997,
28,46,65,91,112,159,361,411,518,612,631,755,895,901,
7,57,75,78,87,224,325,460,494,609,764,800,1028,1034,
31,48,70,79,246,268,437,498,516,572,786,794,1050,1056,
3,34,68,74,110,178,295,448,480,552,626,718,982,988,
30,53,69,78,251,267,436,503,521,571,791,793,1055,1061,
35,38,50,56,72,100,292,308,536,578,591,637,842,848,
18,33,70,89,161,212,321,482,519,673,736,752,1016,1022,
15,24,65,67,175,217,272,278,294,564,604,645,828,834,
36,40,43,66,87,108,300,365,378,648,718,729,912,918,
63,88,89,154,168,260,427,438,453,676,708,769,972,978,
4,58,69,145,164,231,415,473,484,685,748,798,949,955,
47,60,85,130,199,232,384,502,532,751,772,783,1036,1042,
3,13,26,50,57,135,405,486,505,591,675,724,939,945,
9,25,58,61,76,80,331,380,473,594,601,603,865,871,
11,55,73,82,85,222,329,458,492,607,762,798,1026,1032,
4,26,44,79,190,269,357,426,460,595,730,804,994,1000,
19,33,39,81,169,217,396,479,487,707,747,757,1021,1027,
6,21,45,56,234,245,276,374,493,546,683,774,810,816,
9,10,20,146,149,256,329,379,526,561,705,796,1060,1066,
1,55,66,148,167,228,418,470,481,688,745,801,952,958,
11,27,54,63,72,82,333,382,469,596,603,605,867,873,
14,45,74,204,204,223,353,367,474,634,659,744,1008,1014,
3,42,61,119,195,238,297,503,508,609,671,778,1042,1048,
4,35,36,138,142,216,335,389,408,639,654,678,942,948,
6,11,22,145,148,252,325,381,522,563,707,792,1056,1062,
20,30,46,50,53,107,290,292,303,560,743,808,824,830,
14,29,64,66,174,216,271,277,299,569,603,644,833,839,
3,45,87,87,155,160,351,405,430,700,722,773,964,970,
0,31,38,138,140,218,331,385,410,641,656,680,944,950,
9,59,77,80,89,226,327,456,496,611,766,802,1030,1036,
7,12,13,47,183,242,283,311,514,540,553,689,817,823,
20,37,40,55,98,215,368,509,510,551,638,684,902,908,
10,26,59,62,77,81,332,381,468,595,602,604,866,872,
38,50,58,124,167,205,285,437,442,586,707,713,971,977,
42,55,78,89,116,201,282,312,399,582,648,739,846,852,
65,84,85,150,170,262,429,440,455,672,710,771,974,980,
10,16,29,67,99,126,336,396,494,623,664,666,930,936,
64,86,89,199,226,253,314,393,469,571,739,782,1003,1009,
5,15,18,36,61,190,275,358,414,545,564,761,815,1078,
8,13,14,42,184,243,284,306,515,541,554,684,818,824,
2,33,67,73,109,177,294,447,485,557,625,717,981,987,
11,20,44,55,239,244,281,373,492,551,682,779,815,821,
8,17,27,39,57,174,327,345,523,597,650,670,861,867,
23,33,43,50,53,104,289,293,300,563,740,805,827,833,
18,29,76,82,88,137,307,358,375,628,631,696,892,898,
12,27,62,70,178,220,275,281,297,567,601,642,831,837,
25,48,49,65,75,131,319,334,538,580,589,701,853,859,
5,44,63,115,197,234,299,499,504,611,667,774,1038,1044,
7,46,72,92,263,269,365,453,539,561,788,809,1073,1079,
16,47,76,206,206,225,349,369,476,630,655,746,1010,1016,
60,85,88,201,222,255,316,395,471,573,741,784,1005,1011,
30,34,35,55,181,193,300,442,463,569,570,786,834,840,
10,28,77,78,118,210,388,466,524,579,658,763,922,928,
2,44,86,86,154,159,350,404,429,699,721,772,963,969,
4,14,23,41,60,189,274,357,419,544,569,760,814,1077,
6,28,55,64,73,83,334,383,470,597,600,604,868,874,
49,57,69,135,151,256,421,477,487,557,691,713,955,961,
38,40,47,70,85,112,304,363,382,652,716,727,916,922,
10,54,72,81,84,227,328,457,497,606,767,803,1031,1037,
32,49,71,80,247,269,432,499,517,573,787,795,1051,1057,
2,17,73,74,82,191,315,344,461,543,614,626,878,884,
9,15,28,66,98,131,341,401,493,622,663,671,935,941,
30,31,35,56,182,194,301,443,464,564,571,787,835,841,
2,12,21,39,64,187,272,355,417,542,567,758,812,1075,
15,46,75,205,205,224,348,368,475,635,654,745,1009,1015,
7,16,26,38,56,179,326,344,522,596,649,669,860,866,
29,60,67,79,79,250,321,349,412,619,642,663,883,889,
19,34,71,84,156,213,322,483,520,674,737,753,1017,1023,
25,62,69,81,81,246,323,351,408,621,644,665,885,891,
20,36,39,63,123,180,395,423,450,551,720,757,984,990,
24,48,53,64,74,130,318,333,537,579,588,700,852,858,
13,18,19,103,169,239,373,419,531,614,643,777,907,913,
43,56,79,84,117,202,283,313,400,583,649,740,847,853,
23,36,39,60,120,183,392,420,453,548,723,760,987,993,
0,28,46,81,186,265,359,428,456,597,726,806,990,996,
34,37,49,55,77,99,291,307,535,577,590,636,841,847,
8,15,21,52,103,195,275,421,465,719,735,763,999,1005,
5,27,45,80,191,264,358,427,461,596,731,805,995,1001,
9,12,28,40,58,175,328,346,524,598,651,671,862,868,
21,38,41,56,99,210,369,504,511,546,639,685,903,909,
23,31,37,79,173,221,400,477,491,705,745,761,1025,1031,
29,47,60,92,113,160,362,412,519,613,632,750,896,902,
10,11,21,144,147,257,324,380,527,562,706,797,1061,1067,
25,43,62,94,109,156,364,408,521,615,634,752,898,904,
0,15,72,77,80,189,313,342,459,541,612,624,876,882,
32,41,53,59,75,97,289,311,539,581,588,640,845,851,
16,25,60,68,176,218,273,279,295,565,605,646,829,835,
2,56,67,149,162,229,419,471,482,689,746,802,953,959,
0,45,64,116,192,235,294,500,505,606,668,775,1039,1045,
18,37,40,61,121,184,393,421,454,549,724,761,988,994,
4,14,27,51,58,136,406,487,506,592,676,725,940,946,
3,34,41,141,143,221,334,388,413,638,659,683,947,953,
9,13,28,69,249,260,434,445,530,690,694,800,1064,1070,
30,50,63,123,167,228,280,393,446,663,679,792,927,933,
20,34,40,82,170,218,397,474,488,702,748,758,1022,1028,
5,47,89,89,151,156,353,407,426,696,724,769,960,966,
39,41,42,71,86,113,305,364,383,653,717,728,917,923,
34,51,67,82,249,265,434,501,519,575,789,797,1053,1059,
7,13,26,70,96,129,339,399,497,620,661,669,933,939,
1,43,85,85,153,158,349,403,428,698,720,771,962,968,
27,50,51,61,77,127,321,330,534,576,591,697,855,861,
7,22,46,57,235,240,277,375,494,547,678,775,811,817,
8,23,47,58,236,241,278,376,495,548,679,776,812,818,
0,42,84,84,152,157,348,402,427,697,725,770,961,967,
6,13,19,50,107,193,273,425,463,717,733,767,997,1003,
3,4,71,76,78,240,371,404,510,620,731,780,1044,1050,
33,34,35,54,180,192,305,441,462,568,575,791,839,845,
23,32,69,88,160,211,320,481,518,672,735,751,1015,1021,
6,12,17,46,182,241,282,310,513,545,552,688,816,822,
65,84,87,200,227,254,315,394,470,572,740,783,1004,1010,
28,51,52,62,72,128,322,331,535,577,592,698,856,862,
31,32,33,58,184,196,303,439,466,566,573,789,837,843,
13,44,73,209,209,222,352,366,479,633,658,749,1013,1019,
27,45,64,90,111,158,360,410,517,617,630,754,894,900,
37,49,57,123,166,204,284,436,441,585,706,712,970,976,
2,33,40,140,142,220,333,387,412,637,658,682,946,952,
21,26,73,79,85,134,310,355,372,625,634,699,889,895,
6,7,23,146,149,253,326,382,523,558,702,793,1057,1063,
8,9,19,145,148,255,328,378,525,560,704,795,1059,1065,
29,52,53,63,73,129,323,332,536,578,593,699,857,863,
0,5,67,72,80,242,367,406,512,622,727,782,1046,1052,
8,12,27,68,248,259,433,444,529,693,695,799,1063,1069,
2,3,70,75,83,245,370,403,515,619,730,785,1049,1055,
19,35,45,49,52,106,289,291,302,559,742,807,823,829,
44,63,88,127,202,229,387,499,529,754,769,780,1033,1039,
24,61,68,80,80,251,322,350,413,620,643,664,884,890,
45,64,89,128,203,230,388,500,530,755,770,781,1034,1040,
35,49,62,122,166,233,279,392,445,662,678,797,926,932,
0,1,68,73,81,243,368,407,513,623,728,783,1047,1053,
		others => 0);
	end function;

	function init_vector_shifts return vector_shifts is
	begin
		return (
36,18,21,33,46,0,37,45,0,50,7,0,0,0,
0,37,45,9,58,12,0,16,34,0,33,49,0,0,
37,19,21,34,46,0,37,46,0,51,7,0,0,0,
31,15,36,49,34,0,34,46,0,0,19,4,0,0,
33,58,41,49,31,0,32,25,0,54,38,0,0,0,
39,55,0,13,10,0,37,0,32,9,1,0,0,0,
34,58,41,49,31,0,32,25,0,54,38,0,0,0,
0,36,45,58,8,11,0,16,34,0,32,49,0,0,
25,29,31,57,0,17,15,19,0,38,0,30,0,0,
50,39,59,54,52,0,54,0,49,12,31,0,0,0,
53,37,32,19,34,0,30,0,42,5,44,0,0,0,
48,30,42,0,50,8,4,0,24,47,0,31,0,0,
4,42,36,0,47,59,0,31,3,16,54,0,0,0,
33,58,41,48,31,0,32,25,0,54,37,0,0,0,
8,36,20,45,0,12,0,58,55,0,14,45,0,0,
54,47,0,23,5,44,0,53,31,31,0,36,0,0,
16,24,1,11,0,50,0,0,55,0,37,28,0,0,
17,25,1,11,0,51,1,0,55,0,38,29,0,0,
0,8,34,24,27,44,0,29,50,0,31,13,0,0,
9,57,19,0,33,38,23,0,43,0,54,7,0,0,
40,33,31,0,26,56,3,29,0,45,14,0,0,0,
51,39,0,55,53,0,55,0,50,13,32,0,0,0,
13,58,9,37,19,0,49,0,28,18,0,15,0,0,
9,37,20,45,0,13,0,58,56,0,15,46,0,0,
26,26,53,0,27,19,42,0,54,0,43,14,0,0,
33,57,41,48,31,0,32,24,0,53,37,0,0,0,
35,15,0,4,49,2,0,31,6,34,0,5,0,0,
37,43,18,9,0,10,0,4,49,32,0,13,0,0,
37,42,17,8,0,10,0,3,49,32,0,13,0,0,
16,24,1,11,0,50,1,0,55,0,38,28,0,0,
51,39,0,55,53,0,54,0,49,12,32,0,0,0,
0,47,59,53,7,30,0,16,25,0,5,30,0,0,
56,16,36,0,7,38,0,39,4,47,0,51,0,0,
10,47,5,0,6,24,0,27,2,0,11,18,0,0,
6,4,44,44,0,50,55,13,0,21,0,6,0,0,
7,0,26,58,27,10,48,0,37,0,42,49,0,0,
18,6,53,3,0,5,0,3,31,51,0,26,0,0,
56,16,36,0,7,37,0,38,3,47,0,51,0,0,
22,22,26,20,7,0,8,24,0,0,9,18,0,0,
48,31,42,0,50,9,4,0,25,47,0,31,0,0,
26,26,53,0,27,19,42,0,54,0,43,14,0,0,
55,48,38,33,46,0,8,40,0,9,0,37,0,0,
0,13,35,30,33,7,50,0,45,0,27,10,0,0,
18,31,46,47,11,0,56,37,0,35,0,35,0,0,
50,9,17,37,33,0,0,29,49,2,0,16,0,0,
50,54,53,32,43,0,17,8,0,28,5,0,0,0,
13,48,50,31,42,0,5,8,0,18,0,41,0,0,
33,52,11,44,38,0,59,42,0,26,55,0,0,0,
22,22,26,20,6,0,8,24,0,0,9,17,0,0,
33,53,12,45,38,0,59,43,0,26,56,0,0,0,
54,38,47,32,45,0,8,39,0,9,0,36,0,0,
13,48,50,30,42,0,5,8,0,18,0,41,0,0,
50,54,52,32,43,0,17,8,0,5,27,0,0,0,
3,42,35,0,46,58,0,30,2,15,0,53,0,0,
34,28,2,34,0,29,44,0,12,29,0,8,0,0,
30,7,41,47,0,11,29,0,31,30,0,59,0,0,
11,48,5,0,6,24,0,28,3,0,12,19,0,0,
16,24,1,11,0,50,0,0,54,0,37,28,0,0,
33,52,12,44,38,0,59,42,0,26,55,0,0,0,
38,54,59,12,9,0,36,0,31,8,0,0,0,0,
37,42,17,8,0,9,0,3,49,32,0,13,0,0,
39,54,0,13,10,0,36,0,31,9,1,0,0,0,
18,6,52,2,0,4,0,3,31,51,0,26,0,0,
22,21,26,20,6,0,8,24,0,0,8,17,0,0,
18,6,52,2,0,4,0,3,30,50,0,25,0,0,
57,40,38,0,15,32,0,53,14,50,0,14,0,0,
6,4,44,45,0,50,55,13,0,22,0,6,0,0,
54,38,47,32,45,0,8,39,0,9,0,36,0,0,
8,56,19,0,32,37,23,0,42,0,53,6,0,0,
31,8,42,48,0,11,30,0,32,31,0,59,0,0,
25,25,53,0,27,18,41,0,53,0,42,13,0,0,
18,31,46,47,11,0,57,37,0,36,0,35,0,0,
14,59,10,37,20,0,50,0,28,19,0,16,0,0,
31,1,3,29,51,0,8,32,0,58,6,0,0,0,
57,40,38,0,15,32,0,53,14,50,0,14,0,0,
22,4,18,0,52,37,15,55,0,26,0,42,0,0,
33,28,43,24,0,41,0,29,29,46,0,34,0,0,
4,11,7,0,28,32,0,5,51,18,0,22,0,0,
50,9,18,38,33,0,0,29,49,2,0,16,0,0,
0,13,35,30,33,8,50,0,46,0,27,10,0,0,
14,55,0,33,47,9,0,1,15,55,0,4,0,0,
6,0,34,2,28,53,55,13,0,0,57,28,0,0,
51,54,53,33,44,0,17,8,0,28,5,0,0,0,
35,15,0,4,48,2,0,31,6,34,0,5,0,0,
57,40,39,0,16,32,54,0,14,51,0,15,0,0,
0,13,35,30,34,8,50,0,46,0,27,10,0,0,
4,11,7,0,28,32,0,5,52,18,0,23,0,0,
48,31,42,0,51,9,4,0,25,47,0,31,0,0,
18,31,46,48,11,0,57,37,0,36,0,35,0,0,
0,47,59,52,7,30,0,15,25,0,5,30,0,0,
13,58,10,37,20,0,49,0,28,19,0,16,0,0,
51,39,59,54,52,0,54,0,49,12,31,0,0,0,
33,28,43,24,0,41,0,29,29,46,0,34,0,0,
0,37,46,9,58,12,17,0,34,0,33,50,0,0,
4,11,7,0,28,32,0,5,51,18,0,22,0,0,
53,37,32,19,35,0,30,0,43,5,44,0,0,0,
8,57,19,0,32,37,23,0,43,0,53,6,0,0,
0,8,34,24,27,43,0,28,50,0,31,13,0,59,
0,9,34,24,27,44,0,29,50,0,31,13,0,0,
10,47,5,0,6,24,0,28,2,0,11,19,0,0,
23,19,4,0,53,37,15,56,0,26,0,42,0,0,
37,42,17,8,0,9,0,3,49,31,0,12,0,0,
7,0,34,2,28,53,56,14,0,0,57,29,0,0,
33,27,42,23,0,40,0,28,28,45,0,33,0,0,
34,28,2,34,0,29,45,0,12,29,0,9,0,0,
37,43,18,9,0,10,0,4,49,32,0,13,0,0,
52,36,32,19,34,0,30,0,42,5,43,0,0,0,
59,57,28,8,49,0,13,26,0,30,42,0,0,0,
30,7,42,48,0,11,30,0,32,31,0,59,0,0,
57,40,39,0,16,32,54,0,14,51,0,15,0,0,
14,55,0,33,47,9,0,1,15,55,0,4,0,0,
11,33,2,0,51,56,45,18,0,12,39,0,0,0,
50,53,52,32,43,0,17,7,0,27,4,0,0,0,
33,58,41,48,31,0,32,24,0,53,37,0,0,0,
30,7,42,48,0,11,29,0,32,31,0,59,0,0,
48,31,42,0,51,9,5,0,25,48,0,31,0,0,
4,7,10,0,28,31,0,4,51,18,0,22,0,0,
57,40,39,0,16,32,54,0,14,51,0,15,0,0,
41,33,31,27,0,56,3,29,0,46,14,0,0,0,
9,36,20,45,0,12,0,58,55,0,15,45,0,0,
33,2,27,33,0,28,44,0,11,28,0,8,0,0,
34,28,2,34,0,28,44,0,12,29,0,8,0,0,
0,14,35,30,34,8,50,0,46,0,27,11,0,0,
10,33,1,0,51,56,45,18,0,12,39,0,0,0,
8,0,26,58,28,10,48,0,37,0,42,50,0,0,
50,10,18,38,33,0,0,30,50,2,0,17,0,0,
18,6,52,2,0,4,0,3,31,51,0,25,0,0,
31,1,3,29,51,0,9,33,0,59,6,0,0,0,
18,6,52,2,0,4,0,3,30,51,0,25,0,0,
35,15,0,4,49,3,0,31,6,34,0,5,0,0,
9,57,19,0,33,38,24,0,43,0,54,7,0,0,
23,5,19,0,53,37,16,56,0,26,0,43,0,0,
17,31,46,47,10,0,56,36,0,35,0,34,0,0,
31,2,4,30,51,0,9,33,0,59,7,0,0,0,
25,29,31,57,0,17,15,19,0,39,0,31,0,0,
50,10,18,38,33,0,0,29,50,2,0,16,0,0,
33,43,27,24,0,40,0,28,28,45,0,33,0,0,
4,11,7,0,28,32,0,5,52,19,0,23,0,0,
8,0,26,58,28,11,49,0,37,0,42,50,0,0,
57,40,39,0,16,32,54,0,14,50,0,15,0,0,
6,3,43,44,0,50,55,13,0,21,0,6,0,0,
55,15,35,0,6,37,0,38,3,47,0,50,0,0,
13,48,50,31,42,0,5,8,0,18,0,41,0,0,
25,29,30,57,0,16,14,19,0,38,0,30,0,0,
51,39,0,55,53,0,55,0,50,13,32,0,0,0,
26,29,31,58,0,17,15,19,0,39,0,31,0,0,
7,0,26,58,28,10,48,0,37,0,42,50,0,0,
39,54,59,12,9,0,36,0,31,9,0,0,0,0,
6,0,33,2,28,53,55,13,0,0,56,28,0,0,
22,21,26,20,6,0,8,23,0,0,8,17,0,0,
33,27,1,33,0,28,44,0,11,28,0,8,0,0,
10,47,5,0,6,24,0,27,2,0,11,19,0,0,
13,59,10,37,20,0,50,0,28,19,0,16,0,0,
50,10,18,38,33,0,0,30,50,2,0,16,0,0,
3,42,35,0,46,58,0,30,2,16,0,53,0,0,
12,48,50,30,42,0,4,8,0,18,0,41,0,0,
6,4,44,45,0,50,55,14,0,22,0,7,0,0,
31,1,3,29,51,0,9,32,0,58,6,0,0,0,
0,46,58,52,7,29,0,15,25,0,4,30,0,0,
59,57,28,8,49,0,13,27,0,30,42,0,0,0,
11,48,6,0,6,25,0,28,3,0,12,19,0,0,
3,42,36,0,47,58,0,30,3,16,0,53,0,0,
10,32,1,0,51,56,44,18,0,11,38,0,0,0,
33,53,12,44,38,0,59,42,0,26,55,0,0,0,
40,32,31,0,26,56,2,28,0,45,14,0,0,0,
57,58,27,49,7,0,13,26,0,29,41,0,0,0,
0,37,45,58,8,11,0,16,34,0,32,49,0,0,
7,0,34,3,29,54,56,14,0,0,57,29,0,0,
31,15,36,49,33,0,34,46,0,0,19,3,0,0,
41,33,31,27,0,56,3,29,0,45,14,0,0,0,
13,48,50,31,42,0,5,9,0,18,0,41,0,0,
35,15,0,3,48,2,0,30,5,34,0,4,0,0,
33,43,27,24,0,40,0,28,29,45,0,34,0,0,
3,42,35,0,46,58,0,30,3,16,0,53,0,0,
31,8,42,48,0,12,30,0,32,31,0,59,0,0,
0,13,35,29,33,7,50,0,45,0,27,10,0,0,
33,28,2,34,0,28,44,0,11,29,0,8,0,0,
52,36,31,19,34,0,30,0,42,4,43,0,0,0,
22,4,18,0,52,37,15,55,0,26,0,42,0,0,
0,9,35,25,28,44,0,29,51,0,32,13,0,0,
35,15,0,4,48,2,0,31,5,34,0,5,0,0,
51,39,0,55,53,0,55,0,49,12,32,0,0,0,
0,47,59,53,7,30,0,16,26,0,5,30,0,0,
9,36,20,45,0,13,0,58,56,0,15,45,0,0,
0,37,46,9,58,12,17,0,35,0,33,50,0,0,
17,24,1,11,0,50,1,0,55,0,38,29,0,0,
7,0,34,2,28,53,55,13,0,0,57,29,0,0,
54,47,0,22,5,43,0,53,31,31,0,35,0,0,
32,52,11,44,37,0,58,42,0,25,55,0,0,0,
34,58,42,49,31,0,32,25,0,54,38,0,0,0,
10,32,1,0,51,56,45,18,0,12,39,0,0,0,
23,19,4,0,53,37,15,55,0,26,0,42,0,0,
0,13,54,33,47,9,0,0,15,54,0,4,0,0,
18,6,52,3,0,5,0,3,31,51,0,26,0,0,
31,15,36,49,33,0,34,46,0,0,19,3,0,0,
0,9,34,24,28,44,0,29,50,0,31,13,0,0,
4,42,36,0,47,58,0,30,3,16,54,0,0,0,
37,42,17,8,0,9,0,3,49,31,0,12,0,0,
22,22,26,20,7,0,8,24,0,0,9,18,0,0,
13,49,51,31,43,0,5,9,0,19,0,41,0,0,
25,29,30,57,0,16,15,19,0,38,0,30,0,0,
48,30,42,0,50,8,4,0,24,47,0,31,0,0,
53,37,32,20,35,0,30,0,43,5,44,0,0,0,
55,0,13,33,47,9,0,0,15,55,0,4,0,0,
0,9,34,24,27,44,0,29,50,0,31,13,0,0,
10,32,1,0,51,56,45,18,0,11,39,0,0,0,
9,36,20,45,0,12,0,58,56,0,15,45,0,0,
25,26,53,0,27,18,41,0,53,0,43,13,0,0,
39,54,59,13,10,0,36,0,31,9,0,0,0,0,
26,26,53,0,27,19,41,0,54,0,43,13,0,0,
54,38,47,32,45,0,7,39,0,8,0,36,0,0,
54,0,46,22,5,43,0,53,31,31,0,35,0,0,
4,11,7,0,28,31,0,4,51,18,0,22,0,0,
0,13,35,30,33,7,50,0,45,0,27,10,0,0,
54,48,38,33,46,0,8,40,0,9,0,36,0,0,
6,3,43,44,0,50,54,13,0,21,0,6,0,0,
7,0,26,58,27,10,48,0,37,0,42,50,0,0,
18,31,46,47,11,0,56,37,0,35,0,35,0,0,
6,4,44,45,0,51,55,14,0,22,0,7,0,0,
9,37,20,45,0,13,0,58,56,0,15,45,0,0,
33,43,27,24,0,41,0,29,29,46,0,34,0,0,
31,2,4,30,51,0,9,33,0,59,7,0,0,0,
55,15,36,0,6,37,0,38,3,47,0,51,0,0,
59,57,28,50,8,0,14,27,0,30,42,0,0,0,
56,16,36,0,7,38,0,39,3,47,0,51,0,0,
48,30,0,41,50,8,4,0,24,47,0,31,0,0,
8,0,26,58,28,11,49,0,37,0,43,50,0,0,
6,0,34,2,28,53,55,13,0,0,56,28,0,0,
11,48,6,0,7,25,0,28,3,0,12,19,0,0,
33,52,11,44,38,0,59,42,0,26,55,0,0,0,
55,48,38,33,46,0,8,40,0,9,0,36,0,0,
50,10,18,38,33,0,0,30,50,2,0,16,0,0,
41,33,31,27,0,56,3,29,0,46,14,0,0,0,
50,54,52,32,43,0,17,8,0,5,27,0,0,0,
9,57,19,0,32,38,23,0,43,0,54,7,0,0,
31,1,3,29,51,0,9,33,0,59,6,0,0,0,
30,14,35,48,33,0,33,45,0,0,18,3,0,0,
22,22,27,20,7,0,8,24,0,0,9,18,0,0,
25,29,31,57,0,17,15,19,0,38,0,30,0,0,
53,37,32,19,35,0,30,0,42,5,44,0,0,0,
31,15,36,49,33,0,34,46,0,0,19,3,0,0,
54,47,0,23,5,44,0,54,32,32,0,36,0,0,
0,46,58,52,7,30,0,15,25,0,5,30,0,0,
0,46,58,52,7,30,0,15,25,0,5,30,0,0,
31,15,36,49,33,0,34,46,0,0,18,3,0,0,
18,31,46,47,10,0,56,36,0,35,0,34,0,0,
36,18,20,33,46,0,36,45,0,50,6,0,0,0,
14,55,0,34,48,10,0,1,16,55,0,4,0,0,
38,54,59,12,9,0,36,0,31,9,0,0,0,0,
35,0,14,3,48,2,0,30,5,33,0,4,0,0,
22,19,4,0,52,37,15,55,0,26,0,42,0,0,
54,47,0,23,6,44,0,54,32,32,0,36,0,0,
14,55,0,33,47,9,0,1,15,55,0,4,0,0,
11,33,2,0,51,57,45,19,0,12,39,0,0,0,
55,15,35,0,6,37,0,38,3,46,0,50,0,0,
31,8,42,48,0,12,30,0,32,31,0,59,0,0,
41,33,31,27,0,56,3,29,0,46,14,0,0,0,
16,24,1,11,0,50,0,0,55,0,37,28,0,0,
59,57,27,49,7,0,13,26,0,30,42,0,0,0,
59,57,28,8,49,0,13,27,0,30,42,0,0,0,
54,47,0,23,6,44,0,54,32,32,0,36,0,0,
19,36,21,34,46,0,37,45,0,50,7,0,0,0,
50,54,52,32,43,0,17,8,0,27,4,0,0,0,
37,19,21,34,46,0,37,46,0,51,7,0,0,0,
0,36,45,58,8,11,0,16,34,0,32,49,0,0,
13,58,9,37,19,0,49,0,28,18,0,16,0,0,
26,26,53,0,27,18,41,0,53,0,43,13,0,0,
13,58,9,37,19,0,49,0,28,18,0,16,0,0,
8,57,19,0,32,37,23,0,43,0,54,6,0,0,
37,19,21,34,46,0,37,45,0,50,7,0,0,0,
		others => 0);
	end function;
end package body;
