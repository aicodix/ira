-- code table generated from table_vector.txt by generate_table_vector_vhd.cc
--
-- Copyright 2019 Ahmet Inan <inan@aicodix.de>

use work.ldpc_scalar.all;
use work.ldpc_vector.all;

package table_vector is
	function init_vector_parities return vector_parities;
	function init_vector_counts return vector_counts;
	function init_vector_offsets return vector_offsets;
	function init_vector_shifts return vector_shifts;
end package;

package body table_vector is
	function init_vector_parities return vector_parities is
	begin
		return 540;
	end function;

	function init_vector_counts return vector_counts is
	begin
		return (
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
		others => count_scalar'low);
	end function;

	function init_vector_offsets return vector_offsets is
	begin
		return (
8,62,102,134,180,278,672,674,686,1169,1214,1470,1742,1754,
65,103,128,242,328,467,561,782,895,1322,1356,1589,1850,1862,
80,82,95,142,169,226,610,729,766,1306,1430,1459,1834,1846,
94,113,160,177,234,403,574,634,799,1174,1300,1487,1702,1714,
4,85,128,228,394,479,592,996,1019,1222,1338,1559,2087,2099,
23,30,36,103,208,384,542,844,924,1436,1464,1528,1992,2004,
1,29,38,74,129,372,541,714,830,1081,1136,1519,1621,2148,
60,98,123,249,335,462,556,789,890,1329,1363,1584,1857,1869,
49,122,141,159,165,498,647,699,816,1239,1292,1331,1767,1779,
45,61,89,96,105,210,585,587,610,1125,1476,1613,1653,1665,
40,51,152,164,170,267,617,710,751,1250,1271,1396,1778,1790,
11,57,93,158,383,528,712,859,923,1196,1463,1609,1991,2003,
4,5,138,155,157,481,738,813,1021,1239,1458,1561,2089,2101,
35,40,41,215,347,477,755,831,1063,1224,1295,1549,1823,1835,
2,63,76,278,286,442,663,771,826,1279,1318,1366,1894,1906,
30,91,144,412,418,449,705,737,952,1262,1317,1492,2020,2032,
99,119,137,275,309,510,849,953,975,1111,1389,1417,1917,1929,
28,89,154,410,416,447,703,735,950,1260,1315,1490,2018,2030,
20,47,95,118,470,487,560,748,987,1100,1357,1556,1628,1640,
69,107,120,246,332,459,553,786,899,1326,1360,1593,1854,1866,
6,60,100,132,190,276,672,682,684,1167,1212,1468,1740,1752,
49,85,122,184,223,312,724,822,1043,1233,1264,1508,1792,1804,
130,168,179,311,337,519,854,877,910,1349,1417,1538,1945,1957,
89,120,175,256,403,466,774,1006,1066,1501,1546,1569,2074,2086,
14,33,39,106,211,387,545,847,927,1439,1467,1531,1995,2007,
62,77,101,113,147,199,583,617,1079,1157,1182,1276,1685,1697,
4,88,172,178,306,323,706,814,863,1403,1443,1542,1931,1943,
0,34,59,107,114,264,804,981,1018,1176,1344,1441,1872,1884,
60,62,67,117,369,393,602,882,933,1135,1142,1574,1670,1682,
63,101,126,240,326,465,559,780,893,1320,1366,1587,1848,1860,
103,111,141,267,301,514,841,957,979,1115,1381,1421,1909,1921,
91,122,177,258,405,456,776,996,1056,1503,1536,1571,2064,2076,
20,21,37,289,298,507,658,762,1047,1118,1406,1587,2115,2127,
3,64,140,146,218,358,589,898,966,1104,1256,1438,1966,1978,
68,83,107,119,153,193,577,623,1073,1163,1176,1282,1691,1703,
122,171,172,303,341,523,858,881,902,1353,1421,1542,1949,1961,
21,33,52,132,200,257,677,797,991,1246,1323,1337,1865,1877,
13,32,38,105,210,386,544,846,926,1438,1466,1530,1994,2006,
42,53,154,166,172,269,619,712,753,1252,1261,1398,1780,1792,
45,80,83,110,195,426,735,1014,1027,1092,1275,1369,1803,1815,
46,72,81,111,196,427,736,1015,1028,1093,1276,1370,1804,1816,
62,97,143,158,499,539,864,997,1039,1149,1579,1593,2107,2119,
4,31,147,148,162,379,629,688,919,1091,1228,1258,1756,1768,
23,29,34,87,367,486,569,621,1022,1084,1109,1377,1637,1649,
75,77,90,137,176,221,605,724,761,1301,1437,1454,1829,1841,
7,68,81,279,283,435,668,776,819,1272,1311,1359,1887,1899,
37,65,93,97,100,214,577,579,602,1117,1480,1617,1645,1657,
84,115,162,179,236,405,564,624,801,1164,1302,1477,1692,1704,
9,70,134,152,224,352,595,892,960,1110,1250,1432,1960,1972,
64,99,133,160,501,529,866,999,1041,1151,1581,1595,2109,2121,
77,79,92,139,178,223,607,726,763,1303,1439,1456,1831,1843,
14,24,51,134,500,517,871,888,1057,1385,1389,1597,2125,2137,
93,124,179,260,407,458,778,998,1058,1505,1538,1561,2066,2078,
55,91,128,190,217,318,730,816,1037,1227,1270,1502,1798,1810,
13,88,144,188,527,533,725,909,1073,1119,1574,1613,2141,2153,
93,112,159,176,233,402,573,633,798,1173,1299,1486,1701,1713,
11,33,58,106,113,275,815,980,1017,1187,1355,1440,1883,1895,
15,16,44,293,296,514,653,757,1054,1125,1413,1594,2122,2134,
37,70,137,168,318,429,646,969,1036,1346,1475,1509,2037,2049,
129,178,179,310,336,518,853,876,909,1348,1416,1537,1944,1956,
11,60,73,283,287,439,660,768,823,1276,1315,1363,1891,1903,
6,67,80,278,282,434,667,775,818,1283,1310,1358,1886,1898,
19,111,147,162,171,446,655,916,986,1215,1526,1604,2054,2066,
50,98,103,126,154,252,638,671,1079,1163,1178,1392,1706,1718,
13,14,42,291,294,512,651,767,1052,1123,1411,1592,2120,2132,
5,66,79,277,281,433,666,774,817,1282,1309,1357,1885,1897,
85,116,163,168,237,406,565,625,802,1165,1303,1478,1693,1705,
22,29,47,102,207,395,541,843,935,1435,1475,1527,2003,2015,
40,74,83,125,251,362,781,851,902,1099,1442,1515,1970,1982,
8,89,120,232,386,471,596,1000,1011,1214,1342,1551,2079,2091,
42,70,86,102,105,207,582,584,607,1122,1485,1610,1650,1662,
1,115,138,298,335,456,838,944,961,1378,1495,1599,1906,1918,
62,64,69,119,371,395,604,884,935,1137,1144,1576,1672,1684,
70,73,97,109,155,195,579,613,1075,1153,1178,1272,1681,1693,
15,24,58,76,118,349,658,694,1052,1198,1299,1337,1726,1738,
3,87,171,177,305,322,705,813,862,1402,1442,1541,1930,1942,
68,106,131,245,331,458,552,785,898,1325,1359,1592,1853,1865,
1,67,107,139,185,283,677,679,691,1174,1219,1475,1747,1759,
3,84,127,239,393,478,591,1007,1018,1221,1337,1558,2086,2098,
0,27,144,155,158,375,625,684,915,1087,1224,1254,1752,1764,
70,96,121,247,333,460,554,787,888,1327,1361,1594,1855,1867,
128,177,178,309,347,517,852,887,908,1347,1427,1536,1955,1967,
9,31,56,104,111,273,813,978,1015,1185,1353,1450,1881,1893,
57,93,130,180,219,320,720,818,1039,1229,1260,1504,1788,1800,
72,102,116,248,333,413,571,873,884,1166,1413,1419,1941,1953,
20,32,51,143,199,256,676,796,990,1245,1322,1336,1864,1876,
13,35,50,133,499,516,870,899,1056,1384,1388,1596,2124,2136,
36,62,74,158,336,438,803,958,978,1414,1496,1518,2046,2058,
42,68,80,164,342,432,797,952,972,1408,1490,1512,2040,2052,
7,53,89,166,379,536,708,855,919,1192,1459,1617,1987,1999,
18,27,49,79,109,352,649,685,1055,1189,1302,1340,1717,1729,
36,74,83,113,198,429,738,1017,1030,1095,1278,1372,1806,1818,
44,75,78,129,243,366,785,843,906,1103,1446,1519,1974,1986,
87,118,165,170,239,396,567,627,792,1167,1305,1480,1695,1707,
61,99,124,250,324,463,557,790,891,1330,1364,1585,1858,1870,
29,46,47,209,341,471,749,837,1057,1230,1289,1555,1817,1829,
11,92,123,235,389,474,599,1003,1014,1217,1333,1554,2082,2094,
24,85,150,412,418,455,699,743,958,1268,1311,1498,2026,2038,
51,87,124,186,225,314,726,824,1033,1235,1266,1510,1794,1806,
20,112,148,163,172,447,656,917,987,1216,1527,1605,2055,2067,
1,28,144,145,159,376,626,685,916,1088,1225,1255,1753,1765,
70,105,139,166,495,535,872,1005,1035,1145,1575,1589,2103,2115,
79,97,111,243,328,408,566,868,879,1173,1408,1426,1936,1948,
4,32,41,77,120,375,544,717,833,1084,1139,1522,1624,2151,
17,92,148,180,519,537,729,901,1077,1123,1578,1617,2145,2157,
55,128,135,159,165,492,641,705,822,1245,1286,1325,1773,1785,
43,78,81,108,193,424,733,1012,1025,1102,1273,1379,1801,1813,
33,54,125,139,355,433,542,554,594,1134,1210,1293,1662,1674,
18,93,149,181,520,538,730,902,1078,1124,1579,1618,2146,2158,
22,23,39,288,291,509,648,764,1049,1120,1408,1589,2117,2129,
1,62,138,144,216,356,599,896,964,1114,1254,1436,1964,1976,
85,128,171,252,399,462,770,1002,1062,1509,1542,1565,2070,2082,
2,30,39,75,130,373,542,715,831,1082,1137,1520,1622,2149,
14,15,43,292,295,513,652,756,1053,1124,1412,1593,2121,2133,
32,53,124,138,354,432,541,553,593,1133,1209,1292,1661,1673,
54,102,107,130,146,256,642,663,1071,1155,1182,1396,1710,1722,
18,19,47,296,299,505,656,760,1045,1116,1404,1585,2113,2125,
8,69,133,151,223,351,594,891,971,1109,1249,1431,1959,1971,
5,33,42,78,121,376,545,718,834,1085,1128,1523,1625,2152,
4,26,51,99,118,268,808,973,1010,1180,1348,1445,1876,1888,
65,80,104,116,150,202,586,620,1070,1160,1185,1279,1688,1700,
125,171,174,398,449,512,633,790,938,1142,1478,1563,2006,2018,
16,17,45,294,297,515,654,758,1055,1126,1414,1595,2123,2135,
12,52,109,124,151,161,664,761,944,1191,1200,1204,1732,1744,
44,60,88,104,107,209,584,586,609,1124,1487,1612,1652,1664,
54,90,127,189,216,317,729,827,1036,1226,1269,1501,1797,1809,
74,76,89,136,175,220,604,723,760,1300,1436,1453,1828,1840,
123,172,173,304,342,524,859,882,903,1354,1422,1543,1950,1962,
26,87,152,408,414,445,701,733,948,1270,1313,1488,2016,2028,
105,113,143,269,303,504,843,959,981,1105,1383,1423,1911,1923,
47,61,73,157,347,437,802,957,977,1413,1495,1517,2045,2057,
4,70,98,142,188,286,680,682,694,1165,1222,1466,1750,1762,
46,67,134,177,315,426,643,966,1033,1355,1472,1506,2034,2046,
90,109,156,173,230,399,570,630,795,1170,1296,1483,1698,1710,
10,91,122,234,388,473,598,1002,1013,1216,1332,1553,2081,2093,
94,125,168,261,396,459,779,999,1059,1506,1539,1562,2067,2079,
6,52,88,165,378,535,719,854,918,1191,1458,1616,1986,1998,
10,26,47,83,126,381,550,711,839,1090,1133,1516,1630,2157,
0,93,124,236,390,475,588,1004,1015,1218,1334,1555,2083,2095,
37,48,149,161,179,264,614,719,748,1259,1268,1393,1787,1799,
25,86,151,413,419,444,700,732,959,1269,1312,1499,2027,2039,
43,71,87,103,106,208,583,585,608,1123,1486,1611,1651,1663,
7,8,141,146,160,484,741,804,1024,1242,1461,1564,2092,2104,
31,92,145,413,419,450,706,738,953,1263,1318,1493,2021,2033,
16,25,59,77,119,350,659,695,1053,1199,1300,1338,1727,1739,
71,97,122,248,334,461,555,788,889,1328,1362,1595,1856,1868,
17,44,92,115,479,484,557,745,984,1097,1366,1553,1625,1637,
41,69,85,101,104,206,581,583,606,1121,1484,1609,1649,1661,
3,31,40,76,131,374,543,716,832,1083,1138,1521,1623,2150,
18,54,151,164,234,428,774,924,1054,1163,1314,1527,1842,1854,
23,86,154,186,525,531,723,907,1071,1117,1572,1611,2139,2151,
66,104,129,243,329,456,562,783,896,1323,1357,1590,1851,1863,
8,30,55,103,110,272,812,977,1014,1184,1352,1449,1880,1892,
13,25,56,136,192,261,681,801,995,1238,1327,1341,1869,1881,
0,114,137,297,334,467,837,943,960,1377,1494,1598,1905,1917,
72,74,87,134,173,218,602,721,758,1298,1434,1463,1826,1838,
9,55,91,156,381,538,710,857,921,1194,1461,1619,1989,2001,
2,86,170,176,304,321,704,812,861,1401,1441,1540,1929,1941,
8,69,82,280,284,436,669,777,820,1273,1312,1360,1888,1900,
27,48,131,133,349,439,548,560,588,1128,1204,1287,1656,1668,
17,28,35,93,361,480,575,615,1028,1090,1115,1371,1643,1655,
44,65,132,175,313,424,641,964,1043,1353,1470,1504,2032,2044,
6,7,140,145,159,483,740,815,1023,1241,1460,1563,2091,2103,
127,176,177,308,346,516,863,886,907,1346,1426,1547,1954,1966,
72,82,85,132,171,216,600,731,756,1296,1432,1461,1824,1836,
18,24,29,94,362,481,564,616,1029,1091,1104,1372,1632,1644,
7,91,169,175,309,314,697,805,854,1394,1446,1545,1922,1934,
67,105,130,244,330,457,563,784,897,1324,1358,1591,1852,1864,
30,36,47,210,342,472,750,838,1058,1231,1290,1556,1818,1830,
17,53,150,163,233,427,773,935,1053,1162,1313,1526,1841,1853,
86,129,172,253,400,463,771,1003,1063,1510,1543,1566,2071,2083,
5,27,52,100,119,269,809,974,1011,1181,1349,1446,1877,1889,
33,94,147,409,415,452,696,740,955,1265,1308,1495,2023,2035,
35,84,149,411,417,454,698,742,957,1267,1310,1497,2025,2037,
44,55,144,156,174,271,621,714,755,1254,1263,1400,1782,1794,
53,126,133,157,163,502,639,703,820,1243,1284,1323,1771,1783,
86,117,164,169,238,407,566,626,803,1166,1304,1479,1694,1706,
3,64,77,279,287,443,664,772,827,1280,1319,1367,1895,1907,
121,170,179,406,445,508,629,786,946,1150,1486,1571,2014,2026,
40,68,84,100,103,205,580,582,605,1120,1483,1608,1648,1660,
22,50,119,122,149,159,662,759,942,1189,1202,1210,1730,1742,
8,35,151,152,166,383,633,692,923,1083,1232,1250,1760,1772,
78,80,93,140,179,224,608,727,764,1304,1428,1457,1832,1844,
126,175,176,307,345,527,862,885,906,1345,1425,1546,1953,1965,
66,81,105,117,151,203,587,621,1071,1161,1186,1280,1689,1701,
22,34,53,133,201,258,678,798,992,1247,1324,1338,1866,1878,
10,11,132,149,163,487,732,807,1027,1245,1452,1567,2095,2107,
47,63,91,98,107,212,577,587,600,1127,1478,1615,1655,1667,
26,43,44,206,338,468,746,834,1066,1227,1286,1552,1814,1826,
19,25,30,95,363,482,565,617,1030,1080,1105,1373,1633,1645,
10,71,72,282,286,438,671,779,822,1275,1314,1362,1890,1902,
42,73,76,127,241,364,783,841,904,1101,1444,1517,1972,1984,
3,4,137,154,156,480,737,812,1020,1238,1457,1560,2088,2100,
104,112,142,268,302,515,842,958,980,1104,1382,1422,1910,1922,
67,82,106,118,152,192,576,622,1072,1162,1187,1281,1690,1702,
16,56,113,128,155,165,668,765,936,1195,1204,1208,1736,1748,
15,51,148,161,231,425,771,933,1051,1160,1311,1524,1839,1851,
23,38,86,109,473,490,563,751,990,1103,1360,1559,1631,1643,
21,57,154,167,237,431,777,927,1045,1154,1317,1530,1845,1857,
43,74,77,128,242,365,784,842,905,1102,1445,1518,1973,1985,
76,78,91,138,177,222,606,725,762,1302,1438,1455,1830,1842,
34,55,126,140,356,434,543,555,595,1135,1211,1294,1663,1675,
80,98,112,244,329,409,567,869,880,1174,1409,1427,1937,1949,
11,95,173,179,301,318,701,809,858,1398,1450,1537,1926,1938,
41,72,75,126,240,363,782,840,903,1100,1443,1516,1971,1983,
45,71,83,167,345,435,800,955,975,1411,1493,1515,2043,2055,
1,2,135,152,166,490,735,810,1030,1236,1455,1570,2098,2110,
61,76,100,112,146,198,582,616,1078,1156,1181,1275,1684,1696,
71,74,98,110,144,196,580,614,1076,1154,1179,1273,1682,1694,
11,26,154,155,157,374,624,695,914,1086,1235,1253,1763,1775,
10,94,172,178,300,317,700,808,857,1397,1449,1536,1925,1937,
12,48,145,158,228,422,768,930,1048,1157,1308,1533,1836,1848,
38,71,138,169,319,430,647,970,1037,1347,1464,1510,2038,2050,
1,62,75,277,285,441,662,770,825,1278,1317,1365,1893,1905,
12,13,41,290,293,511,650,766,1051,1122,1410,1591,2119,2131,
10,56,92,157,382,539,711,858,922,1195,1462,1608,1990,2002,
69,104,138,165,494,534,871,1004,1034,1144,1574,1588,2102,2114,
12,39,87,110,474,491,552,752,991,1092,1361,1548,1620,1632,
0,84,168,174,302,319,702,810,859,1399,1451,1538,1927,1939,
20,56,153,166,236,430,776,926,1044,1153,1316,1529,1844,1856,
3,69,97,141,187,285,679,681,693,1164,1221,1465,1749,1761,
87,130,173,254,401,464,772,1004,1064,1511,1544,1567,2072,2084,
15,90,146,190,517,535,727,911,1075,1121,1576,1615,2143,2155,
11,60,136,154,226,354,597,894,962,1112,1252,1434,1962,1974,
6,108,143,291,328,461,831,937,966,1371,1488,1604,1899,1911,
73,103,117,249,334,414,572,874,885,1167,1414,1420,1942,1954,
20,30,57,140,494,523,865,894,1063,1383,1391,1603,2131,2143,
13,49,146,159,229,423,769,931,1049,1158,1309,1534,1837,1849,
52,125,132,156,162,501,638,702,819,1242,1295,1322,1770,1782,
57,130,137,161,167,494,643,707,824,1247,1288,1327,1775,1787,
59,120,139,157,163,496,645,697,826,1237,1290,1329,1765,1777,
107,115,133,271,305,506,845,949,983,1107,1385,1425,1913,1925,
20,27,45,100,205,393,551,841,933,1433,1473,1525,2001,2013,
35,56,127,141,357,435,544,556,596,1136,1200,1295,1664,1676,
0,1,134,151,165,489,734,809,1029,1247,1454,1569,2097,2109,
17,26,48,78,108,351,648,684,1054,1188,1301,1339,1716,1728,
16,27,34,92,360,491,574,614,1027,1089,1114,1370,1642,1654,
43,64,143,174,312,423,640,963,1042,1352,1469,1503,2031,2043,
5,32,148,149,163,380,630,689,920,1080,1229,1259,1757,1769,
2,95,126,238,392,477,590,1006,1017,1220,1336,1557,2085,2097,
40,75,78,117,202,421,742,1009,1022,1099,1282,1376,1810,1822,
64,69,71,114,366,390,611,879,930,1132,1151,1583,1679,1691,
2,63,139,145,217,357,588,897,965,1115,1255,1437,1965,1977,
39,67,95,99,102,204,579,581,604,1119,1482,1619,1647,1659,
28,45,46,208,340,470,748,836,1056,1229,1288,1554,1816,1828,
47,68,135,178,316,427,644,967,1034,1344,1473,1507,2035,2047,
1,59,95,160,373,530,714,861,913,1198,1453,1611,1981,1993,
8,110,133,293,330,463,833,939,968,1373,1490,1606,1901,1913,
41,76,79,118,203,422,743,1010,1023,1100,1283,1377,1811,1823,
1,35,48,96,115,265,805,982,1019,1177,1345,1442,1873,1885,
88,119,166,171,228,397,568,628,793,1168,1306,1481,1696,1708,
12,116,152,167,176,451,648,921,991,1220,1531,1597,2059,2071,
78,96,110,242,327,419,565,867,878,1172,1407,1425,1935,1947,
9,25,46,82,125,380,549,710,838,1089,1132,1515,1629,2156,
40,61,140,171,321,420,637,960,1039,1349,1466,1500,2028,2040,
84,127,170,263,398,461,769,1001,1061,1508,1541,1564,2069,2081,
65,100,134,161,502,530,867,1000,1042,1140,1582,1584,2110,2122,
16,28,59,139,195,252,672,792,986,1241,1330,1332,1860,1872,
31,52,123,137,353,443,540,552,592,1132,1208,1291,1660,1672,
9,10,143,148,162,486,743,806,1026,1244,1463,1566,2094,2106,
4,118,141,289,326,459,829,947,964,1369,1498,1602,1897,1909,
1,85,169,175,303,320,703,811,860,1400,1440,1539,1928,1940,
3,117,140,288,325,458,828,946,963,1368,1497,1601,1896,1908,
6,87,130,230,384,469,594,998,1009,1212,1340,1549,2077,2089,
79,81,94,141,168,225,609,728,765,1305,1429,1458,1833,1845,
15,25,52,135,501,518,872,889,1058,1386,1390,1598,2126,2138,
16,43,91,114,478,483,556,744,995,1096,1365,1552,1624,1636,
21,31,58,141,495,524,866,895,1064,1380,1384,1604,2132,2144,
81,99,113,245,330,410,568,870,881,1175,1410,1416,1938,1950,
2,3,136,153,167,491,736,811,1031,1237,1456,1571,2099,2111,
17,18,46,295,298,504,655,759,1044,1127,1415,1584,2112,2124,
22,31,53,83,113,356,653,689,1047,1193,1306,1332,1721,1733,
124,173,174,305,343,525,860,883,904,1355,1423,1544,1951,1963,
19,94,150,182,521,539,731,903,1079,1125,1580,1619,2147,2159,
50,86,123,185,224,313,725,823,1032,1234,1265,1509,1793,1805,
21,36,84,119,471,488,561,749,988,1101,1358,1557,1629,1641,
19,46,94,117,469,486,559,747,986,1099,1356,1555,1627,1639,
15,42,90,113,477,482,555,755,994,1095,1364,1551,1623,1635,
81,83,84,143,170,227,611,730,767,1307,1431,1460,1835,1847,
31,36,37,211,343,473,751,839,1059,1232,1291,1557,1819,1831,
10,71,135,153,225,353,596,893,961,1111,1251,1433,1961,1973,
39,73,82,124,250,361,780,850,901,1098,1441,1514,1969,1981,
8,92,170,176,310,315,698,806,855,1395,1447,1546,1923,1935,
46,62,90,97,106,211,576,586,611,1126,1477,1614,1654,1666,
19,55,152,165,235,429,775,925,1055,1152,1315,1528,1843,1855,
131,168,169,300,338,520,855,878,911,1350,1418,1539,1946,1958,
56,129,136,160,166,493,642,706,823,1246,1287,1326,1774,1786,
5,119,142,290,327,460,830,936,965,1370,1499,1603,1898,1910,
16,108,144,159,168,455,652,913,995,1212,1535,1601,2063,2075,
44,70,82,166,344,434,799,954,974,1410,1492,1514,2042,2054,
48,96,101,124,152,262,636,669,1077,1161,1176,1402,1704,1716,
63,98,132,159,500,528,865,998,1040,1150,1580,1594,2108,2120,
42,77,80,119,192,423,732,1011,1024,1101,1272,1378,1800,1812,
50,123,142,160,166,499,636,700,817,1240,1293,1320,1768,1780,
17,29,48,140,196,253,673,793,987,1242,1331,1333,1861,1873,
56,97,104,120,148,258,644,665,1073,1157,1184,1398,1712,1724,
37,72,75,114,199,430,739,1018,1031,1096,1279,1373,1807,1819,
19,59,116,131,146,156,671,756,939,1198,1207,1211,1739,1751,
67,102,136,163,492,532,869,1002,1032,1142,1572,1586,2100,2112,
9,70,83,281,285,437,670,778,821,1274,1313,1361,1889,1901,
95,114,161,178,235,404,575,635,800,1175,1301,1476,1703,1715,
51,99,104,127,155,253,639,660,1068,1152,1179,1393,1707,1719,
130,176,179,403,454,505,626,783,943,1147,1483,1568,2011,2023,
6,34,43,79,122,377,546,719,835,1086,1129,1512,1626,2153,
54,127,134,158,164,503,640,704,821,1244,1285,1324,1772,1784,
41,52,153,165,171,268,618,711,752,1251,1260,1397,1779,1791,
3,25,50,98,117,267,807,972,1009,1179,1347,1444,1875,1887,
60,107,141,156,497,537,874,1007,1037,1147,1577,1591,2105,2117,
43,69,81,165,343,433,798,953,973,1409,1491,1513,2041,2053,
82,100,114,246,331,411,569,871,882,1164,1411,1417,1939,1951,
124,170,173,397,448,511,632,789,937,1141,1477,1562,2005,2017,
129,175,178,402,453,504,625,782,942,1146,1482,1567,2010,2022,
0,61,74,276,284,440,661,769,824,1277,1316,1364,1892,1904,
4,65,141,147,219,359,590,899,967,1105,1257,1439,1967,1979,
1,94,125,237,391,476,589,1005,1016,1219,1335,1556,2084,2096,
45,66,133,176,314,425,642,965,1032,1354,1471,1505,2033,2045,
74,104,118,250,335,415,573,875,886,1168,1415,1421,1943,1955,
101,109,139,265,311,512,851,955,977,1113,1391,1419,1919,1931,
120,169,178,405,444,507,628,785,945,1149,1485,1570,2013,2025,
14,26,57,137,193,262,682,802,984,1239,1328,1342,1870,1882,
7,61,101,133,191,277,673,683,685,1168,1213,1469,1741,1753,
5,66,142,148,220,348,591,888,968,1106,1258,1428,1956,1968,
123,169,172,396,447,510,631,788,936,1140,1476,1561,2004,2016,
38,73,76,115,200,431,740,1019,1020,1097,1280,1374,1808,1820,
128,174,177,401,452,515,624,781,941,1145,1481,1566,2009,2021,
58,94,131,181,220,321,721,819,1040,1230,1261,1505,1789,1801,
106,114,132,270,304,505,844,948,982,1106,1384,1424,1912,1924,
24,57,128,142,358,436,545,557,597,1137,1201,1284,1665,1677,
83,101,115,247,332,412,570,872,883,1165,1412,1418,1940,1952,
25,58,129,143,359,437,546,558,598,1138,1202,1285,1666,1678,
73,75,88,135,174,219,603,722,759,1299,1435,1452,1827,1839,
12,23,40,289,292,510,649,765,1050,1121,1409,1590,2118,2130,
0,11,133,150,164,488,733,808,1028,1246,1453,1568,2096,2108,
2,48,84,161,374,531,715,862,914,1199,1454,1612,1982,1994,
28,49,120,134,350,440,549,561,589,1129,1205,1288,1657,1669,
63,65,70,108,360,384,605,885,924,1138,1145,1577,1673,1685,
22,85,153,185,524,530,722,906,1070,1116,1583,1610,2138,2150,
18,30,49,141,197,254,674,794,988,1243,1320,1334,1862,1874,
5,71,99,143,189,287,681,683,695,1166,1223,1467,1751,1763,
32,93,146,408,414,451,707,739,954,1264,1319,1494,2022,2034,
2,68,96,140,186,284,678,680,692,1175,1220,1464,1748,1760,
37,80,83,122,248,371,790,848,911,1096,1451,1512,1979,1991,
76,106,108,240,325,417,575,865,876,1170,1405,1423,1933,1945,
36,59,148,160,178,275,613,718,747,1258,1267,1392,1786,1798,
66,101,135,162,503,531,868,1001,1043,1141,1583,1585,2111,2123,
61,96,142,157,498,538,875,996,1038,1148,1578,1592,2106,2118,
89,108,167,172,229,398,569,629,794,1169,1307,1482,1697,1709,
59,100,107,123,151,261,647,668,1076,1160,1187,1401,1715,1727,
20,48,117,120,147,157,660,757,940,1199,1200,1208,1728,1740,
23,32,54,72,114,357,654,690,1048,1194,1307,1333,1722,1734,
38,66,94,98,101,215,578,580,603,1118,1481,1618,1646,1658,
19,26,44,99,204,392,550,840,932,1432,1472,1524,2000,2012,
56,92,129,191,218,319,731,817,1038,1228,1271,1503,1799,1811,
62,67,69,112,364,388,609,877,928,1130,1149,1581,1677,1689,
48,121,140,158,164,497,646,698,827,1238,1291,1330,1766,1778,
96,116,134,272,306,507,846,950,972,1108,1386,1426,1914,1926,
51,124,143,161,167,500,637,701,818,1241,1294,1321,1769,1781,
97,117,135,273,307,508,847,951,973,1109,1387,1427,1915,1927,
45,76,79,130,244,367,786,844,907,1092,1447,1520,1975,1987,
4,50,86,163,376,533,717,852,916,1189,1456,1614,1984,1996,
37,63,75,159,337,439,792,959,979,1415,1497,1519,2047,2059,
47,78,81,120,246,369,788,846,909,1094,1449,1522,1977,1989,
16,91,147,191,518,536,728,900,1076,1122,1577,1616,2144,2156,
126,172,175,399,450,513,634,791,939,1143,1479,1564,2007,2019,
69,72,96,108,154,194,578,612,1074,1152,1177,1283,1680,1692,
19,20,36,288,297,506,657,761,1046,1117,1405,1586,2114,2126,
16,26,53,136,502,519,873,890,1059,1387,1391,1599,2127,2139,
13,40,88,111,475,480,553,753,992,1093,1362,1549,1621,1633,
7,29,54,102,109,271,811,976,1013,1183,1351,1448,1879,1891,
0,61,137,155,227,355,598,895,963,1113,1253,1435,1963,1975,
3,49,85,162,375,532,716,863,915,1188,1455,1613,1983,1995,
13,117,153,156,177,452,649,922,992,1221,1532,1598,2060,2072,
60,75,99,111,145,197,581,615,1077,1155,1180,1274,1683,1695,
23,33,48,143,497,526,868,897,1066,1382,1386,1606,2134,2146,
19,31,50,142,198,255,675,795,989,1244,1321,1335,1863,1875,
7,34,150,151,165,382,632,691,922,1082,1231,1249,1759,1771,
0,66,106,138,184,282,676,678,690,1173,1218,1474,1746,1758,
20,29,51,81,111,354,651,687,1045,1191,1304,1342,1719,1731,
12,33,55,73,115,358,655,691,1049,1195,1296,1334,1723,1735,
36,79,82,121,247,370,789,847,910,1095,1450,1523,1978,1990,
38,72,81,123,249,360,791,849,900,1097,1440,1513,1968,1980,
20,26,31,84,364,483,566,618,1031,1081,1106,1374,1634,1646,
14,35,57,75,117,348,657,693,1051,1197,1298,1336,1725,1737,
5,89,173,179,307,312,707,815,852,1392,1444,1543,1920,1932,
21,22,38,290,299,508,659,763,1048,1119,1407,1588,2116,2128,
46,77,80,131,245,368,787,845,908,1093,1448,1521,1976,1988,
61,66,68,111,363,387,608,876,927,1129,1148,1580,1676,1688,
47,58,147,159,177,274,612,717,746,1257,1266,1403,1785,1797,
7,109,132,292,329,462,832,938,967,1372,1489,1605,1900,1912,
39,50,151,163,169,266,616,709,750,1249,1270,1395,1777,1789,
63,68,70,113,365,389,610,878,929,1131,1150,1582,1678,1690,
125,174,175,306,344,526,861,884,905,1344,1424,1545,1952,1964,
14,54,111,126,153,163,666,763,946,1193,1202,1206,1734,1746,
39,65,77,161,339,441,794,949,981,1405,1499,1521,2049,2061,
18,45,93,116,468,485,558,746,985,1098,1367,1554,1626,1638,
17,109,145,160,169,444,653,914,984,1213,1524,1602,2052,2064,
46,60,72,156,346,436,801,956,976,1412,1494,1516,2044,2056,
15,119,155,158,179,454,651,912,994,1223,1534,1600,2062,2074,
13,24,31,89,369,488,571,623,1024,1086,1111,1379,1639,1651,
18,58,115,130,145,167,670,767,938,1197,1206,1210,1738,1750,
10,64,104,136,182,280,674,676,688,1171,1216,1472,1744,1756,
102,110,140,266,300,513,840,956,978,1114,1380,1420,1908,1920,
7,88,131,231,385,470,595,999,1010,1213,1341,1550,2078,2090,
21,84,152,184,523,529,721,905,1069,1127,1582,1609,2137,2149,
62,100,125,251,325,464,558,791,892,1331,1365,1586,1859,1871,
68,103,137,164,493,533,870,1003,1033,1143,1573,1587,2101,2113,
33,38,39,213,345,475,753,829,1061,1234,1293,1559,1821,1833,
27,88,153,409,415,446,702,734,949,1271,1314,1489,2017,2029,
11,113,136,296,333,466,836,942,971,1376,1493,1597,1904,1916,
34,39,40,214,346,476,754,830,1062,1235,1294,1548,1822,1834,
64,79,103,115,149,201,585,619,1069,1159,1184,1278,1687,1699,
98,118,136,274,308,509,848,952,974,1110,1388,1416,1916,1928,
10,112,135,295,332,465,835,941,970,1375,1492,1596,1903,1915,
42,63,142,173,323,422,639,962,1041,1351,1468,1502,2030,2042,
57,98,105,121,149,259,645,666,1074,1158,1185,1399,1713,1725,
12,30,35,88,368,487,570,622,1023,1085,1110,1378,1638,1650,
19,29,56,139,493,522,864,893,1062,1382,1390,1602,2130,2142,
34,95,148,410,416,453,697,741,956,1266,1309,1496,2024,2036,
23,115,151,166,175,450,659,920,990,1219,1530,1596,2058,2070,
21,113,149,164,173,448,657,918,988,1217,1528,1606,2056,2068,
15,34,40,107,212,388,546,848,928,1428,1468,1532,1996,2008,
41,67,79,163,341,443,796,951,983,1407,1489,1523,2051,2063,
92,111,158,175,232,401,572,632,797,1172,1298,1485,1700,1712,
77,107,109,241,326,418,564,866,877,1171,1406,1424,1934,1946,
7,35,44,80,123,378,547,708,836,1087,1130,1513,1627,2154,
9,111,134,294,331,464,834,940,969,1374,1491,1607,1902,1914,
18,25,43,98,215,391,549,851,931,1431,1471,1535,1999,2011,
59,95,120,182,221,322,722,820,1041,1231,1262,1506,1790,1802,
38,49,150,162,168,265,615,708,749,1248,1269,1394,1776,1788,
12,87,155,187,526,532,724,908,1072,1118,1573,1612,2140,2152,
73,83,86,133,172,217,601,720,757,1297,1433,1462,1825,1837,
0,58,94,159,372,529,713,860,912,1197,1452,1610,1980,1992,
10,25,153,154,156,373,635,694,913,1085,1234,1252,1762,1774,
36,64,92,96,99,213,576,578,601,1116,1479,1616,1644,1656,
24,41,42,204,336,478,744,832,1064,1225,1284,1550,1812,1824,
9,63,103,135,181,279,673,675,687,1170,1215,1471,1743,1755,
18,28,55,138,492,521,875,892,1061,1381,1389,1601,2129,2141,
32,37,38,212,344,474,752,828,1060,1233,1292,1558,1820,1832,
75,105,119,251,324,416,574,864,887,1169,1404,1422,1932,1944,
5,86,129,229,395,468,593,997,1008,1223,1339,1548,2076,2088,
29,50,121,135,351,441,550,562,590,1130,1206,1289,1658,1670,
21,30,52,82,112,355,652,688,1046,1192,1305,1343,1720,1732,
20,95,151,183,522,528,720,904,1068,1126,1581,1608,2136,2148,
40,66,78,162,340,442,795,950,982,1406,1488,1522,2050,2062,
52,88,125,187,226,315,727,825,1034,1224,1267,1511,1795,1807,
60,65,70,115,367,391,600,880,931,1133,1140,1572,1668,1680,
120,169,170,301,339,521,856,879,900,1351,1419,1540,1947,1959,
39,74,77,116,201,420,741,1008,1021,1098,1281,1375,1809,1821,
0,28,37,73,128,383,540,713,829,1080,1135,1518,1620,2159,
12,24,55,135,203,260,680,800,994,1237,1326,1340,1868,1880,
49,97,102,125,153,263,637,670,1078,1162,1177,1403,1705,1717,
22,114,150,165,174,449,658,919,989,1218,1529,1607,2057,2069,
9,90,121,233,387,472,597,1001,1012,1215,1343,1552,2080,2092,
30,51,122,136,352,442,551,563,591,1131,1207,1290,1659,1671,
12,34,49,132,498,527,869,898,1067,1383,1387,1607,2135,2147,
53,89,126,188,227,316,728,826,1035,1225,1268,1500,1796,1808,
23,51,108,123,150,160,663,760,943,1190,1203,1211,1731,1743,
91,110,157,174,231,400,571,631,796,1171,1297,1484,1699,1711,
48,84,121,183,222,323,723,821,1042,1232,1263,1507,1791,1803,
2,29,145,146,160,377,627,686,917,1089,1226,1256,1754,1766,
4,65,78,276,280,432,665,773,816,1281,1308,1356,1884,1896,
61,66,71,116,368,392,601,881,932,1134,1141,1573,1669,1681,
64,102,127,241,327,466,560,781,894,1321,1367,1588,1849,1861,
8,54,90,167,380,537,709,856,920,1193,1460,1618,1988,2000,
46,57,146,158,176,273,623,716,745,1256,1265,1402,1784,1796,
6,33,149,150,164,381,631,690,921,1081,1230,1248,1758,1770,
131,168,177,404,455,506,627,784,944,1148,1484,1569,2012,2024,
53,101,106,129,145,255,641,662,1070,1154,1181,1395,1709,1721,
18,110,146,161,170,445,654,915,985,1214,1525,1603,2053,2065,
13,34,56,74,116,359,656,692,1050,1196,1297,1335,1724,1736,
64,66,71,109,361,385,606,886,925,1139,1146,1578,1674,1686,
88,131,174,255,402,465,773,1005,1065,1500,1545,1568,2073,2085,
23,35,54,134,202,259,679,799,993,1236,1325,1339,1867,1879,
21,49,118,121,148,158,661,758,941,1188,1201,1209,1729,1741,
58,99,106,122,150,260,646,667,1075,1159,1186,1400,1714,1726,
45,56,145,157,175,272,622,715,744,1255,1264,1401,1783,1795,
21,27,32,85,365,484,567,619,1020,1082,1107,1375,1635,1647,
127,173,176,400,451,514,635,780,940,1144,1480,1565,2008,2020,
60,65,67,110,362,386,607,887,926,1128,1147,1579,1675,1687,
14,118,154,157,178,453,650,923,993,1222,1533,1599,2061,2073,
15,26,33,91,371,490,573,613,1026,1088,1113,1369,1641,1653,
17,57,114,129,144,166,669,766,937,1196,1205,1209,1737,1749,
14,50,147,160,230,424,770,932,1050,1159,1310,1535,1838,1850,
15,55,112,127,154,164,667,764,947,1194,1203,1207,1735,1747,
8,24,45,81,124,379,548,709,837,1088,1131,1514,1628,2155,
121,170,171,302,340,522,857,880,901,1352,1420,1541,1948,1960,
22,32,59,142,496,525,867,896,1065,1381,1385,1605,2133,2145,
9,24,152,153,167,372,634,693,912,1084,1233,1251,1761,1773,
11,65,105,137,183,281,675,677,689,1172,1217,1473,1745,1757,
47,73,82,112,197,428,737,1016,1029,1094,1277,1371,1805,1817,
17,24,42,97,214,390,548,850,930,1430,1470,1534,1998,2010,
41,62,141,172,322,421,638,961,1040,1350,1467,1501,2029,2041,
122,168,171,407,446,509,630,787,947,1151,1487,1560,2015,2027,
36,69,136,179,317,428,645,968,1035,1345,1474,1508,2036,2048,
3,30,146,147,161,378,628,687,918,1090,1227,1257,1755,1767,
2,116,139,299,324,457,839,945,962,1379,1496,1600,1907,1919,
43,54,155,167,173,270,620,713,754,1253,1262,1399,1781,1793,
63,78,102,114,148,200,584,618,1068,1158,1183,1277,1686,1698,
23,59,144,157,239,421,779,929,1047,1156,1319,1532,1847,1859,
5,51,87,164,377,534,718,853,917,1190,1457,1615,1985,1997,
22,37,85,108,472,489,562,750,989,1102,1359,1558,1630,1642,
44,79,82,109,194,425,734,1013,1026,1103,1274,1368,1802,1814,
29,90,155,411,417,448,704,736,951,1261,1316,1491,2019,2031,
71,106,140,167,496,536,873,1006,1036,1146,1576,1590,2104,2116,
95,126,169,262,397,460,768,1000,1060,1507,1540,1563,2068,2080,
6,28,53,101,108,270,810,975,1012,1182,1350,1447,1878,1890,
61,63,68,118,370,394,603,883,934,1136,1143,1575,1671,1683,
8,9,142,147,161,485,742,805,1025,1243,1462,1565,2093,2105,
16,35,41,96,213,389,547,849,929,1429,1469,1533,1997,2009,
92,123,178,259,406,457,777,997,1057,1504,1537,1560,2065,2077,
15,27,58,138,194,263,683,803,985,1240,1329,1343,1871,1883,
6,90,168,174,308,313,696,804,853,1393,1445,1544,1921,1933,
13,53,110,125,152,162,665,762,945,1192,1201,1205,1733,1745,
22,28,33,86,366,485,568,620,1021,1083,1108,1376,1636,1648,
6,67,143,149,221,349,592,889,969,1107,1259,1429,1957,1969,
90,121,176,257,404,467,775,1007,1067,1502,1547,1570,2075,2087,
19,28,50,80,110,353,650,686,1044,1190,1303,1341,1718,1730,
12,31,37,104,209,385,543,845,925,1437,1465,1529,1993,2005,
100,108,138,264,310,511,850,954,976,1112,1390,1418,1918,1930,
21,28,46,101,206,394,540,842,934,1434,1474,1526,2002,2014,
10,32,57,105,112,274,814,979,1016,1186,1354,1451,1882,1894,
14,89,145,189,516,534,726,910,1074,1120,1575,1614,2142,2154,
39,60,139,170,320,431,636,971,1038,1348,1465,1511,2039,2051,
25,42,43,205,337,479,745,833,1065,1226,1285,1551,1813,1825,
58,131,138,156,162,495,644,696,825,1236,1289,1328,1764,1776,
5,6,139,144,158,482,739,814,1022,1240,1459,1562,2090,2102,
38,64,76,160,338,440,793,948,980,1404,1498,1520,2048,2060,
17,27,54,137,503,520,874,891,1060,1380,1388,1600,2128,2140,
52,100,105,128,144,254,640,661,1069,1153,1180,1394,1708,1720,
22,58,155,156,238,420,778,928,1046,1155,1318,1531,1846,1858,
27,44,45,207,339,469,747,835,1067,1228,1287,1553,1815,1827,
14,25,32,90,370,489,572,612,1025,1087,1112,1368,1640,1652,
16,52,149,162,232,426,772,934,1052,1161,1312,1525,1840,1852,
7,68,132,150,222,350,593,890,970,1108,1248,1430,1958,1970,
9,93,171,177,311,316,699,807,856,1396,1448,1547,1924,1936,
14,41,89,112,476,481,554,754,993,1094,1363,1550,1622,1634,
55,96,103,131,147,257,643,664,1072,1156,1183,1397,1711,1723,
11,27,36,72,127,382,551,712,828,1091,1134,1517,1631,2158,
26,59,130,132,348,438,547,559,599,1139,1203,1286,1667,1679,
2,24,49,97,116,266,806,983,1008,1178,1346,1443,1874,1886,
		others => 0);
	end function;

	function init_vector_shifts return vector_shifts is
	begin
		return (
28,20,19,0,8,16,27,0,7,25,0,7,0,0,
4,28,9,0,16,18,11,0,21,0,27,3,0,0,
11,11,13,10,4,0,4,12,0,0,5,9,0,0,
0,7,18,15,17,4,25,0,23,0,14,5,0,0,
17,27,6,23,19,0,0,22,0,13,28,0,0,0,
8,15,23,23,5,0,28,18,0,17,0,17,0,0,
0,4,17,12,13,22,0,14,25,0,15,6,0,0,
5,29,10,0,16,19,12,0,22,0,27,4,0,0,
13,13,26,0,13,9,20,0,27,0,21,6,0,0,
0,19,23,5,29,6,0,8,17,0,17,25,0,0,
8,12,0,5,0,25,0,0,27,0,18,14,0,0,
3,2,22,23,0,26,28,7,0,11,0,4,0,0,
18,9,10,16,23,0,18,22,0,25,3,0,0,0,
2,6,4,0,14,16,0,3,26,10,0,12,0,0,
21,17,16,14,0,28,2,15,0,23,7,0,0,0,
5,16,1,0,25,28,22,9,0,6,19,0,0,0,
19,21,9,4,0,5,0,2,25,16,0,7,0,0,
5,16,0,0,25,28,22,9,0,6,19,0,0,0,
0,23,29,26,4,15,0,8,13,0,3,15,0,0,
4,28,10,0,16,19,12,0,21,0,27,3,0,0,
28,20,19,0,7,16,0,26,7,25,0,7,0,0,
28,8,18,0,3,19,0,19,1,23,0,25,0,0,
16,1,13,16,0,14,22,0,5,14,0,4,0,0,
7,0,5,19,10,0,25,0,14,10,0,8,0,0,
9,15,23,23,5,0,28,18,0,17,0,17,0,0,
4,0,13,29,14,5,24,0,18,0,21,25,0,0,
16,8,25,18,17,0,17,23,0,0,10,2,0,0,
25,4,8,18,16,0,0,14,24,1,0,8,0,0,
7,0,27,16,23,4,0,0,7,27,0,2,0,0,
4,28,9,0,16,18,11,0,21,0,26,3,0,0,
18,21,8,4,0,4,0,1,24,15,0,6,0,0,
6,29,4,18,9,0,24,0,14,9,0,7,0,0,
29,28,14,4,24,0,6,13,0,15,21,0,0,0,
26,20,0,28,27,0,28,0,25,7,16,0,0,0,
4,0,13,29,14,6,25,0,19,0,22,25,0,0,
17,14,1,17,0,14,22,0,6,14,0,4,0,0,
26,18,16,10,17,0,15,0,21,2,22,0,0,0,
9,15,23,23,5,0,28,18,0,17,0,17,0,0,
8,12,0,5,0,25,0,0,27,0,19,14,0,0,
16,21,13,12,0,20,0,14,14,23,0,17,0,0,
16,14,21,12,0,20,0,14,14,23,0,17,0,0,
13,15,15,29,0,8,8,10,0,19,0,15,0,0,
24,15,21,0,25,4,2,0,12,23,0,15,0,0,
17,0,7,2,24,1,0,15,3,17,0,2,0,0,
11,11,13,10,3,0,4,12,0,0,4,9,0,0,
20,16,15,0,13,28,1,14,0,23,7,0,0,0,
0,18,22,29,4,5,0,8,17,0,16,24,0,0,
0,6,17,14,16,3,25,0,22,0,13,5,0,0,
25,19,0,27,26,0,27,0,25,6,16,0,0,0,
13,15,16,29,0,9,8,10,0,19,0,15,0,0,
11,11,13,10,3,0,4,12,0,0,4,9,0,0,
25,27,26,16,21,0,8,4,0,2,13,0,0,0,
6,29,4,18,9,0,24,0,14,9,0,8,0,0,
28,8,18,0,4,19,0,20,2,24,0,26,0,0,
17,29,21,24,15,0,16,12,0,27,19,0,0,0,
0,7,18,15,17,4,25,0,23,0,14,5,0,0,
25,5,9,19,17,0,0,15,25,1,0,9,0,0,
0,29,14,25,4,0,7,14,0,15,21,0,0,0,
20,27,0,7,5,0,18,0,16,5,0,0,0,0,
16,13,0,16,0,14,22,0,5,14,0,4,0,0,
20,17,16,0,13,28,2,15,0,23,7,0,0,0,
20,16,15,0,13,28,1,14,0,22,7,0,0,0,
6,24,25,15,21,0,2,4,0,9,0,20,0,0,
27,0,23,11,2,22,0,26,15,15,0,18,0,0,
0,29,14,25,4,0,7,13,0,15,21,0,0,0,
20,16,15,0,13,28,1,14,0,22,7,0,0,0,
0,6,17,15,16,3,25,0,22,0,13,5,0,0,
9,16,23,24,6,0,29,19,0,18,0,18,0,0,
27,19,23,16,22,0,4,19,0,4,0,18,0,0,
16,26,6,22,19,0,29,21,0,13,27,0,0,0,
0,18,23,29,4,6,0,8,17,0,16,25,0,0,
6,24,3,0,3,13,0,14,2,0,6,10,0,0,
7,0,27,16,23,4,0,0,7,27,0,2,0,0,
3,0,13,29,13,5,24,0,18,0,21,25,0,0,
5,19,10,23,0,7,0,29,28,0,8,23,0,0,
16,8,25,18,17,0,17,23,0,0,10,2,0,0,
4,28,9,0,16,19,12,0,21,0,27,3,0,0,
29,20,19,0,8,16,27,0,7,25,0,7,0,0,
17,27,6,22,19,0,0,21,0,13,28,0,0,0,
24,15,0,20,25,4,2,0,12,23,0,15,0,0,
4,29,10,0,16,19,12,0,22,0,27,3,0,0,
17,14,1,17,0,15,23,0,6,15,0,5,0,0,
25,5,9,19,17,0,0,15,25,1,0,8,0,0,
27,7,17,0,3,18,0,19,1,23,0,25,0,0,
16,4,21,24,0,6,15,0,16,16,0,0,0,0,
26,18,16,9,17,0,15,0,21,2,22,0,0,0,
25,26,26,16,21,0,8,3,0,2,13,0,0,0,
16,1,2,15,26,0,4,16,0,29,3,0,0,0,
15,0,1,14,25,0,4,16,0,29,3,0,0,0,
3,2,22,22,0,25,28,7,0,11,0,3,0,0,
4,18,10,22,0,6,0,29,27,0,7,22,0,0,
17,14,21,12,0,20,0,14,14,23,0,17,0,0,
27,24,19,16,23,0,4,20,0,4,0,18,0,0,
0,6,17,15,16,4,25,0,23,0,13,5,0,0,
5,29,10,0,17,19,12,0,22,0,27,4,0,0,
2,5,3,0,14,16,0,2,26,9,0,11,0,0,
16,26,6,22,19,0,29,21,0,13,28,0,0,0,
6,17,1,26,0,28,23,9,0,6,20,0,0,0,
28,8,18,0,3,19,0,19,2,23,0,25,0,0,
6,24,25,15,21,0,2,4,0,9,0,20,0,0,
24,15,21,0,25,4,2,0,12,23,0,15,0,0,
12,14,15,28,0,8,7,9,0,19,0,15,0,0,
15,4,21,24,0,6,15,0,16,15,0,29,0,0,
0,4,17,12,14,22,0,14,25,0,15,6,0,0,
17,29,21,25,16,0,16,13,0,27,19,0,0,0,
13,13,27,14,0,10,21,0,27,0,22,7,0,0,
16,21,13,12,0,20,0,14,14,22,0,16,0,0,
3,0,17,1,14,27,28,7,0,0,28,14,0,0,
17,29,21,25,16,0,16,13,0,27,19,0,0,0,
29,28,14,25,4,0,7,13,0,15,21,0,0,0,
26,20,0,28,27,0,27,0,25,6,16,0,0,0,
7,29,5,19,10,0,25,0,14,9,0,8,0,0,
0,4,17,12,13,22,0,14,25,0,15,6,0,0,
0,29,14,25,4,0,7,14,0,15,21,0,0,0,
3,0,17,1,14,27,28,7,0,0,28,14,0,0,
27,0,23,11,3,22,0,27,16,16,0,18,0,0,
29,28,13,24,3,0,6,13,0,15,21,0,0,0,
25,19,0,27,26,0,27,0,24,6,16,0,0,0,
0,4,17,12,14,22,0,14,25,0,16,6,0,0,
25,5,9,19,16,0,0,15,25,1,0,8,0,0,
4,0,13,29,14,5,24,0,19,0,21,25,0,0,
11,2,9,0,26,18,7,27,0,13,0,21,0,0,
0,29,14,25,4,0,7,14,0,15,21,0,0,0,
2,21,18,0,23,29,0,15,1,8,27,0,0,0,
0,19,23,29,4,6,0,8,17,0,16,25,0,0,
28,8,18,0,4,19,0,19,2,24,0,26,0,0,
11,11,13,10,3,0,4,12,0,0,4,9,0,0,
17,14,1,17,0,14,22,0,6,14,0,4,0,0,
5,16,0,0,25,28,22,9,0,5,19,0,0,0,
18,21,8,4,0,5,0,1,24,16,0,6,0,0,
15,1,2,15,25,0,4,16,0,29,3,0,0,0,
29,20,20,0,8,16,27,0,7,26,0,8,0,0,
19,27,0,6,5,0,18,0,16,4,0,0,0,0,
0,7,18,15,17,4,25,0,23,0,14,5,0,0,
16,26,6,22,19,0,29,21,0,13,28,0,0,0,
6,29,5,18,10,0,24,0,14,9,0,8,0,0,
3,2,22,22,0,25,27,7,0,11,0,3,0,0,
0,5,17,12,14,22,0,15,25,0,16,7,0,0,
17,26,6,22,19,0,0,21,0,13,28,0,0,0,
9,13,1,6,0,26,1,0,28,0,19,15,0,0,
6,17,1,26,0,29,23,10,0,6,20,0,0,0,
0,18,23,29,4,6,0,8,17,0,16,25,0,0,
18,9,10,17,23,0,18,23,0,25,3,0,0,0,
5,16,1,0,25,28,22,9,0,6,19,0,0,0,
5,19,10,23,0,7,0,29,28,0,8,23,0,0,
4,29,10,0,16,19,12,0,22,0,27,3,0,0,
0,23,29,26,3,15,0,8,13,0,2,15,0,0,
0,18,23,29,4,6,0,8,17,0,16,25,0,0,
0,4,17,12,13,22,0,14,25,0,15,6,0,0,
9,3,26,1,0,2,0,2,15,25,0,13,0,0,
16,29,20,24,15,0,16,12,0,27,19,0,0,0,
4,28,9,0,16,19,11,0,21,0,27,3,0,0,
25,5,9,19,17,0,0,15,25,1,0,8,0,0,
27,19,16,10,18,0,15,0,21,3,22,0,0,0,
6,24,3,0,3,12,0,14,2,0,6,10,0,0,
11,11,13,10,3,0,4,12,0,0,4,8,0,0,
3,2,22,23,0,25,28,7,0,11,0,3,0,0,
16,8,25,18,17,0,17,23,0,0,10,2,0,0,
20,16,15,0,13,28,1,14,0,23,7,0,0,0,
3,0,16,1,14,26,27,6,0,0,28,14,0,0,
18,8,0,2,25,2,0,16,3,17,0,3,0,0,
19,27,0,6,5,0,18,0,15,4,0,0,0,0,
18,9,10,17,23,0,18,22,0,25,3,0,0,0,
17,14,1,17,0,15,22,0,6,15,0,4,0,0,
11,10,13,10,3,0,4,11,0,0,4,8,0,0,
17,0,7,1,24,1,0,15,2,16,0,2,0,0,
15,7,18,24,16,0,17,23,0,0,9,1,0,0,
4,28,9,0,16,19,11,0,21,0,27,3,0,0,
2,4,5,0,14,16,0,2,26,9,0,11,0,0,
9,3,26,1,0,2,0,1,15,25,0,13,0,0,
7,29,5,19,10,0,25,0,14,9,0,8,0,0,
25,5,9,19,16,0,0,15,25,1,0,8,0,0,
5,16,1,26,0,28,23,9,0,6,20,0,0,0,
5,17,1,26,0,28,23,9,0,6,20,0,0,0,
8,12,1,6,0,25,0,0,27,0,19,14,0,0,
13,13,27,14,0,9,21,0,27,0,22,7,0,0,
0,6,17,15,16,3,25,0,22,0,13,5,0,0,
21,17,16,14,0,28,2,15,0,23,7,0,0,0,
12,10,2,0,27,19,8,28,0,13,0,21,0,0,
0,18,23,29,4,6,0,8,17,0,16,25,0,0,
1,21,17,0,23,29,0,15,1,8,0,26,0,0,
24,15,21,0,25,4,2,0,12,24,0,16,0,0,
11,11,13,10,3,0,4,12,0,0,5,9,0,0,
17,14,1,17,0,14,22,0,6,15,0,4,0,0,
4,0,13,29,14,5,24,0,19,0,21,25,0,0,
26,18,16,10,17,0,15,0,21,2,22,0,0,0,
18,9,11,17,23,0,19,23,0,25,4,0,0,0,
0,19,23,5,29,6,9,0,18,0,17,25,0,0,
2,5,3,0,14,16,0,2,25,9,0,11,0,0,
17,0,7,1,24,1,0,15,2,17,0,2,0,0,
20,16,16,0,13,28,1,14,0,23,7,0,0,0,
27,24,19,16,23,0,4,20,0,4,0,18,0,0,
18,9,10,16,23,0,18,22,0,25,3,0,0,0,
18,21,8,4,0,4,0,1,24,16,0,6,0,0,
4,0,13,29,14,6,25,0,19,0,21,25,0,0,
2,21,18,0,23,29,0,15,2,8,27,0,0,0,
9,3,26,1,0,2,0,1,15,25,0,13,0,0,
0,24,0,27,4,15,0,8,13,0,3,15,0,0,
9,3,26,1,0,2,0,2,16,26,0,13,0,0,
27,24,19,16,23,0,4,20,0,4,0,18,0,0,
11,11,13,10,3,0,4,12,0,0,4,9,0,0,
3,0,17,1,14,27,28,7,0,0,28,14,0,0,
15,4,21,24,0,6,15,0,16,15,0,29,0,0,
15,7,18,24,17,0,17,23,0,0,9,2,0,0,
27,24,19,16,23,0,4,20,0,4,0,18,0,0,
15,0,1,14,25,0,4,16,0,29,3,0,0,0,
19,10,11,17,23,0,19,23,0,26,4,0,0,0,
4,0,13,29,14,5,24,0,18,0,21,25,0,0,
3,0,13,29,14,5,24,0,18,0,21,25,0,0,
24,16,21,0,26,5,3,0,13,24,0,16,0,0,
15,7,18,24,17,0,17,23,0,0,9,2,0,0,
9,3,26,1,0,2,0,1,15,25,0,12,0,0,
20,27,0,7,5,0,18,0,16,5,1,0,0,0,
21,17,16,14,0,28,2,15,0,23,7,0,0,0,
0,29,14,25,4,0,7,13,0,15,21,0,0,0,
3,2,22,23,0,25,28,7,0,11,0,4,0,0,
12,14,15,28,0,8,7,9,0,19,0,15,0,0,
0,23,29,26,3,14,0,7,12,0,2,15,0,0,
16,8,25,18,17,0,17,23,0,0,9,2,0,0,
9,3,26,1,0,2,0,2,16,26,0,13,0,0,
29,20,20,0,8,16,27,0,7,26,0,8,0,0,
7,29,5,19,10,0,25,0,14,9,0,8,0,0,
17,29,21,24,16,0,16,12,0,27,19,0,0,0,
25,20,0,27,26,0,27,0,25,6,16,0,0,0,
5,24,2,0,3,12,0,14,1,0,6,9,0,0,
16,4,21,24,0,6,15,0,16,16,0,0,0,0,
25,27,26,16,22,0,9,4,0,14,2,0,0,0,
9,3,26,1,0,2,0,1,15,25,0,12,0,0,
13,13,27,14,0,9,21,0,27,0,21,7,0,0,
13,13,27,14,0,10,21,0,27,0,22,7,0,0,
12,13,26,0,13,9,20,0,26,0,21,6,0,0,
18,21,9,4,0,5,0,2,24,16,0,6,0,0,
9,16,23,24,6,0,28,19,0,18,0,18,0,0,
3,0,17,1,14,27,28,7,0,0,29,14,0,0,
19,10,11,17,23,0,19,23,0,25,4,0,0,0,
4,18,10,22,0,6,0,29,27,0,7,22,0,0,
18,8,0,2,25,1,0,16,3,17,0,3,0,0,
19,27,29,6,5,0,18,0,15,4,0,0,0,0,
24,15,21,0,25,4,2,0,12,24,0,15,0,0,
17,26,6,22,19,0,0,21,0,13,28,0,0,0,
17,22,14,12,0,21,0,15,15,23,0,17,0,0,
28,7,0,17,24,5,0,1,8,28,0,2,0,0,
26,20,0,28,27,0,28,0,25,6,16,0,0,0,
0,18,22,29,4,6,0,8,17,0,16,24,0,0,
2,5,3,0,14,16,0,2,26,9,0,11,0,0,
19,27,0,6,5,0,18,0,16,5,0,0,0,0,
3,1,21,22,0,25,27,6,0,10,0,3,0,0,
5,24,3,0,3,12,0,14,1,0,6,9,0,0,
17,22,14,12,0,21,0,15,15,23,0,17,0,0,
25,4,9,19,16,0,0,14,24,1,0,8,0,0,
0,6,17,15,17,4,25,0,23,0,13,5,0,0,
7,24,25,15,21,0,3,4,0,9,0,21,0,0,
15,4,21,24,0,5,15,0,16,15,0,29,0,0,
0,5,17,12,14,22,0,15,25,0,16,7,0,0,
19,27,29,6,4,0,18,0,15,4,0,0,0,0,
7,29,5,18,10,0,25,0,14,9,0,8,0,0,
13,15,16,29,0,9,8,10,0,20,0,16,0,0,
26,18,15,9,17,0,15,0,21,2,21,0,0,0,
3,0,17,1,14,26,28,7,0,0,28,14,0,0,
18,9,10,17,23,0,18,23,0,25,3,0,0,0,
5,23,2,0,3,12,0,13,1,0,5,9,0,0,
16,8,25,18,17,0,17,23,0,0,10,2,0,0,
5,23,2,0,3,12,0,13,1,0,5,9,0,0,
16,26,5,22,19,0,29,21,0,13,27,0,0,0,
11,11,13,10,4,0,4,12,0,0,5,9,0,0,
25,27,26,16,21,0,8,4,0,2,13,0,0,0,
0,23,29,26,3,15,0,8,12,0,2,15,0,0,
25,27,26,16,22,0,9,4,0,3,14,0,0,0,
15,4,21,24,0,6,15,0,16,15,0,0,0,0,
19,10,11,17,23,0,19,23,0,26,4,0,0,0,
29,28,13,24,3,0,6,13,0,14,20,0,0,0,
4,18,10,22,0,6,0,29,28,0,7,23,0,0,
17,14,1,17,0,14,22,0,6,14,0,4,0,0,
17,29,21,25,16,0,16,13,0,27,19,0,0,0,
28,8,18,0,3,19,0,19,2,23,0,25,0,0,
0,24,0,26,4,15,0,8,13,0,3,15,0,0,
0,23,29,26,4,15,0,8,13,0,3,15,0,0,
0,23,29,26,3,15,0,7,12,0,2,15,0,0,
11,11,14,10,4,0,4,12,0,0,5,9,0,0,
2,6,4,0,14,16,0,2,26,9,0,11,0,0,
25,19,0,27,26,0,27,0,25,6,16,0,0,0,
27,19,23,16,22,0,4,19,0,4,0,18,0,0,
15,7,18,24,16,0,17,23,0,0,9,1,0,0,
0,19,23,5,29,6,9,0,17,0,17,25,0,0,
9,3,26,1,0,2,0,2,15,26,0,13,0,0,
16,14,1,17,0,14,22,0,5,14,0,4,0,0,
13,13,27,14,0,10,21,0,27,0,22,7,0,0,
5,23,2,0,3,12,0,14,1,0,5,9,0,0,
7,25,26,16,22,0,3,5,0,10,0,21,0,0,
15,0,1,14,25,0,4,16,0,29,3,0,0,0,
27,0,23,11,2,21,0,26,15,15,0,17,0,0,
13,15,16,29,0,9,8,10,0,19,0,15,0,0,
16,21,13,11,0,20,0,14,14,22,0,16,0,0,
13,13,26,0,13,9,21,0,27,0,21,7,0,0,
26,18,16,9,17,0,15,0,21,2,21,0,0,0,
27,24,0,12,3,22,0,27,16,16,0,18,0,0,
17,22,14,12,0,20,0,14,14,23,0,17,0,0,
2,21,18,0,24,0,0,16,2,8,27,0,0,0,
12,14,15,28,0,8,7,9,0,19,0,15,0,0,
20,16,15,0,13,28,1,14,0,23,7,0,0,0,
0,7,18,15,17,4,25,0,23,0,14,6,0,0,
27,0,23,11,2,22,0,27,16,16,0,18,0,0,
11,2,9,0,26,19,8,28,0,13,0,21,0,0,
0,4,17,12,14,22,0,14,25,0,16,7,0,0,
13,13,27,14,0,9,21,0,27,0,22,7,0,0,
8,12,0,5,0,25,0,0,27,0,19,14,0,0,
25,5,9,19,16,0,0,15,25,1,0,8,0,0,
13,14,15,29,0,8,7,9,0,19,0,15,0,0,
15,0,1,14,25,0,4,16,0,29,3,0,0,0,
15,4,21,24,0,6,15,0,16,16,0,0,0,0,
11,2,9,0,26,18,7,27,0,13,0,21,0,0,
11,2,9,0,26,19,8,28,0,13,0,21,0,0,
21,17,16,14,0,28,2,15,0,23,7,0,0,0,
26,20,0,28,27,0,28,0,25,7,16,0,0,0,
17,26,6,22,19,0,0,21,0,13,28,0,0,0,
19,27,0,6,5,0,18,0,16,4,0,0,0,0,
16,4,21,24,0,6,15,0,16,16,0,0,0,0,
19,22,9,5,0,5,0,2,25,16,0,7,0,0,
12,10,2,0,27,19,8,28,0,13,0,21,0,0,
27,19,16,10,18,0,15,0,22,3,22,0,0,0,
28,20,19,0,7,16,0,26,7,25,0,7,0,0,
25,19,29,27,26,0,27,0,24,6,15,0,0,0,
11,2,9,0,26,18,7,27,0,13,0,21,0,0,
17,22,14,12,0,20,0,14,15,23,0,17,0,0,
11,2,9,0,26,18,8,28,0,13,0,21,0,0,
27,7,17,0,3,18,0,19,1,23,0,25,0,0,
18,21,9,4,0,5,0,2,24,16,0,6,0,0,
4,0,17,1,14,27,28,7,0,0,29,15,0,0,
15,4,21,24,0,6,15,0,16,16,0,0,0,0,
4,0,17,1,14,27,28,7,0,0,29,15,0,0,
11,11,13,10,3,0,4,12,0,0,4,9,0,0,
29,29,14,25,4,0,7,13,0,15,21,0,0,0,
10,18,11,17,23,0,19,23,0,25,4,0,0,0,
3,2,22,22,0,25,27,6,0,10,0,3,0,0,
3,0,17,1,14,26,27,6,0,0,28,14,0,0,
7,0,27,17,24,5,0,0,8,27,0,2,0,0,
16,29,20,24,15,0,16,12,0,27,18,0,0,0,
26,18,16,9,17,0,15,0,21,2,22,0,0,0,
29,20,20,0,8,16,27,0,7,26,0,8,0,0,
5,16,1,26,0,28,22,9,0,6,19,0,0,0,
29,20,20,0,8,16,27,0,7,25,0,8,0,0,
28,24,19,17,23,0,4,20,0,5,0,19,0,0,
15,3,21,24,0,5,14,0,16,15,0,29,0,0,
9,12,1,6,0,25,1,0,28,0,19,15,0,0,
13,15,16,29,0,9,8,10,0,20,0,16,0,0,
13,15,15,29,0,8,7,10,0,19,0,15,0,0,
0,7,17,15,17,4,25,0,23,0,13,5,0,0,
27,24,0,12,3,22,0,27,16,16,0,18,0,0,
1,21,17,0,23,29,0,15,1,7,0,26,0,0,
4,18,10,23,0,6,0,29,28,0,7,23,0,0,
0,18,22,29,4,5,0,8,17,0,16,24,0,0,
9,16,23,24,6,0,28,19,0,18,0,18,0,0,
28,8,18,0,4,19,0,20,2,24,0,26,0,0,
28,7,0,17,24,5,0,1,8,28,0,2,0,0,
13,13,26,0,13,9,20,0,26,0,21,6,0,0,
19,21,9,4,0,5,0,2,25,16,0,6,0,0,
13,13,26,0,13,9,21,0,27,0,21,7,0,0,
19,21,9,4,0,5,0,2,25,16,0,6,0,0,
27,24,19,16,23,0,4,20,0,5,0,18,0,0,
3,2,22,22,0,25,27,7,0,11,0,3,0,0,
16,1,2,15,26,0,5,16,0,29,3,0,0,0,
27,24,19,17,23,0,4,20,0,5,0,18,0,0,
17,29,21,24,16,0,16,13,0,27,19,0,0,0,
11,2,9,0,26,18,7,27,0,13,0,21,0,0,
3,0,13,29,13,5,24,0,18,0,21,24,0,0,
29,28,14,4,24,0,6,13,0,15,21,0,0,0,
25,27,26,16,21,0,8,4,0,2,13,0,0,0,
0,23,29,26,3,15,0,7,12,0,2,15,0,0,
25,5,9,19,17,0,0,15,25,1,0,8,0,0,
26,20,0,27,26,0,27,0,25,6,16,0,0,0,
3,2,22,22,0,25,27,6,0,11,0,3,0,0,
7,24,25,16,21,0,3,4,0,9,0,21,0,0,
4,0,13,29,14,5,24,0,18,0,21,25,0,0,
25,27,27,16,22,0,9,4,0,3,14,0,0,0,
26,18,16,9,17,0,15,0,21,2,22,0,0,0,
24,15,21,0,25,4,2,0,12,24,0,16,0,0,
29,20,19,0,8,16,27,0,7,25,0,7,0,0,
4,18,10,22,0,6,0,29,28,0,7,22,0,0,
5,18,10,23,0,6,0,29,28,0,8,23,0,0,
28,24,19,17,23,0,4,20,0,5,0,18,0,0,
27,19,23,16,22,0,3,19,0,4,0,18,0,0,
17,0,7,2,24,1,0,15,2,17,0,2,0,0,
5,18,10,23,0,7,0,29,28,0,8,23,0,0,
15,7,24,17,16,0,16,22,0,0,9,1,0,0,
29,28,14,4,24,0,6,13,0,15,21,0,0,0,
27,24,19,16,23,0,4,20,0,5,0,18,0,0,
28,7,0,17,24,5,0,1,8,28,0,2,0,0,
8,12,1,6,0,25,1,0,28,0,19,14,0,0,
5,24,3,0,3,12,0,14,1,0,6,9,0,0,
8,12,0,5,0,25,0,0,27,0,18,14,0,0,
28,7,0,17,24,5,0,1,8,28,0,2,0,0,
17,14,1,17,0,14,22,0,6,15,0,4,0,0,
2,21,18,0,23,29,0,15,1,8,27,0,0,0,
16,1,2,15,26,0,5,17,0,0,3,0,0,0,
0,23,29,26,4,15,0,8,13,0,2,15,0,0,
6,24,25,15,21,0,2,4,0,9,0,20,0,0,
15,1,2,15,25,0,4,16,0,29,3,0,0,0,
7,24,25,16,21,0,3,5,0,9,0,21,0,0,
18,8,0,2,24,1,0,15,3,17,0,2,0,0,
2,21,18,0,24,29,0,15,2,8,27,0,0,0,
28,20,19,0,8,16,27,0,7,25,0,7,0,0,
18,21,8,4,0,4,0,1,24,15,0,6,0,0,
16,26,5,22,19,0,29,21,0,13,27,0,0,0,
16,29,20,24,15,0,16,12,0,26,18,0,0,0,
5,29,10,0,17,19,12,0,22,0,27,4,0,0,
12,14,15,28,0,8,7,9,0,19,0,15,0,0,
2,6,4,0,14,16,0,3,26,9,0,11,0,0,
5,16,0,0,25,28,22,9,0,5,19,0,0,0,
5,24,3,0,3,12,0,14,1,0,6,10,0,0,
2,6,4,0,14,16,0,3,26,9,0,12,0,0,
4,0,13,29,14,5,24,0,19,0,21,25,0,0,
19,21,9,4,0,5,0,2,25,16,0,7,0,0,
5,24,3,0,3,12,0,14,1,0,6,10,0,0,
19,27,29,6,4,0,18,0,15,4,0,0,0,0,
27,24,0,12,3,22,0,27,16,16,0,18,0,0,
18,0,7,2,24,1,0,15,3,17,0,2,0,0,
25,27,26,16,22,0,9,4,0,14,2,0,0,0,
5,16,1,26,0,28,23,9,0,6,20,0,0,0,
6,24,25,15,21,0,2,4,0,9,0,21,0,0,
6,24,25,15,21,0,2,4,0,9,0,20,0,0,
9,15,23,23,5,0,28,18,0,18,0,17,0,0,
16,1,2,15,26,0,5,17,0,0,4,0,0,0,
0,7,18,15,17,4,25,0,23,0,14,5,0,0,
15,3,21,24,0,5,15,0,16,15,0,29,0,0,
0,4,17,12,14,22,0,15,25,0,16,7,0,0,
5,24,3,0,3,12,0,14,1,0,6,9,0,0,
9,16,23,24,5,0,28,18,0,18,0,17,0,0,
27,7,18,0,3,18,0,19,1,23,0,25,0,0,
8,12,0,5,0,25,0,0,27,0,18,14,0,0,
17,29,20,24,15,0,16,12,0,27,19,0,0,0,
11,10,13,10,3,0,4,12,0,0,4,8,0,0,
3,1,21,22,0,25,27,6,0,10,0,3,0,0,
24,16,21,0,26,5,2,0,13,24,0,16,0,0,
0,18,22,29,4,5,0,8,17,0,16,24,0,0,
2,5,3,0,14,15,0,2,25,9,0,11,0,0,
28,20,19,0,8,16,27,0,7,25,0,7,0,0,
25,27,26,16,22,0,8,4,0,14,2,0,0,0,
2,6,4,0,14,16,0,3,26,9,0,11,0,0,
15,3,20,23,0,5,14,0,15,15,0,29,0,0,
16,26,5,22,18,0,29,21,0,12,27,0,0,0,
3,0,17,1,14,26,27,6,0,0,28,14,0,0,
4,18,10,22,0,6,0,29,28,0,7,22,0,0,
16,28,20,24,15,0,16,12,0,26,18,0,0,0,
16,1,2,15,26,0,5,17,0,0,4,0,0,0,
28,8,18,0,3,19,0,19,2,24,0,25,0,0,
0,27,6,16,23,4,0,0,7,27,0,2,0,0,
17,14,1,17,0,14,22,0,6,14,0,4,0,0,
17,22,14,12,0,21,0,15,15,23,0,17,0,0,
0,4,17,12,13,21,0,14,25,0,15,6,0,29,
27,19,16,10,17,0,15,0,21,3,22,0,0,0,
27,0,23,11,2,21,0,26,15,15,0,17,0,0,
6,24,25,15,21,0,2,4,0,9,0,20,0,0,
16,26,6,22,19,0,29,21,0,13,27,0,0,0,
3,0,17,1,14,26,27,6,0,0,28,14,0,0,
26,27,27,17,22,0,9,4,0,3,14,0,0,0,
28,8,18,0,3,19,0,19,2,24,0,26,0,0,
1,21,18,0,23,29,0,15,1,8,0,26,0,0,
0,7,18,15,17,4,25,0,23,0,14,5,0,0,
28,8,18,0,3,18,0,19,1,23,0,25,0,0,
24,15,21,0,25,4,2,0,12,23,0,15,0,0,
20,16,15,0,13,28,1,14,0,22,7,0,0,0,
0,27,6,16,23,4,0,0,7,27,0,2,0,0,
4,28,9,0,16,18,11,0,21,0,26,3,0,0,
3,2,22,22,0,25,28,7,0,11,0,3,0,0,
8,12,1,6,0,25,0,0,28,0,19,14,0,0,
24,15,21,0,25,4,2,0,12,24,0,16,0,0,
11,10,2,0,26,19,8,28,0,13,0,21,0,0,
27,0,23,11,3,22,0,27,16,16,0,18,0,0,
6,24,25,15,21,0,2,4,0,9,0,20,0,0,
5,18,10,23,0,6,0,29,28,0,8,23,0,0,
7,0,27,17,24,5,0,0,8,27,0,2,0,0,
7,29,5,19,10,0,25,0,14,10,0,8,0,0,
26,18,16,10,17,0,15,0,21,3,22,0,0,0,
1,21,17,0,23,29,0,15,1,8,0,26,0,0,
27,24,0,12,3,22,0,27,16,16,0,18,0,0,
8,12,1,6,0,25,0,0,28,0,19,14,0,0,
17,0,7,2,24,1,0,15,3,17,0,2,0,0,
11,2,9,0,26,18,7,28,0,13,0,21,0,0,
28,7,0,17,24,5,0,0,8,28,0,2,0,0,
7,24,25,16,21,0,3,4,0,9,0,21,0,0,
18,8,0,2,24,1,0,16,3,17,0,3,0,0,
2,21,18,0,24,29,0,15,2,8,27,0,0,0,
9,3,26,1,0,2,0,1,15,25,0,12,0,0,
2,21,18,0,23,29,0,15,1,8,27,0,0,0,
0,5,17,12,14,22,0,15,25,0,16,7,0,0,
17,14,1,17,0,14,22,0,6,14,0,4,0,0,
25,27,26,16,22,0,9,4,0,3,14,0,0,0,
24,16,21,0,25,5,2,0,13,24,0,16,0,0,
28,20,19,0,8,16,27,0,7,25,0,7,0,0,
16,14,21,12,0,20,0,14,14,23,0,17,0,0,
9,16,23,24,5,0,28,18,0,18,0,17,0,0,
19,27,29,6,4,0,18,0,15,4,0,0,0,0,
12,3,10,0,27,19,8,28,0,13,0,22,0,0,
20,27,0,6,5,0,18,0,16,5,0,0,0,0,
24,15,21,0,25,4,2,0,12,23,0,15,0,0,
6,24,3,0,4,13,0,14,2,0,6,10,0,0,
8,12,0,5,0,25,0,0,27,0,19,14,0,0,
4,0,13,29,14,5,24,0,19,0,21,25,0,0,
9,3,27,2,0,3,0,2,16,26,0,13,0,0,
3,2,22,22,0,25,27,7,0,11,0,3,0,0,
0,24,0,27,4,15,0,8,13,0,3,15,0,0,
16,21,13,12,0,20,0,14,14,22,0,17,0,0,
5,16,0,0,25,28,22,9,0,6,19,0,0,0,
12,14,15,28,0,8,7,9,0,19,0,15,0,0,
6,29,5,18,10,0,25,0,14,9,0,8,0,0,
25,5,9,19,17,0,0,15,25,1,0,8,0,0,
7,0,27,16,23,4,0,0,7,27,0,2,0,0,
18,9,10,17,23,0,18,23,0,25,3,0,0,0,
9,15,23,24,5,0,28,18,0,18,0,17,0,0,
6,29,4,18,9,0,24,0,14,9,0,8,0,0,
27,19,16,10,18,0,15,0,22,3,22,0,0,0,
15,7,18,24,16,0,17,23,0,0,9,1,0,0,
2,21,18,0,23,29,0,15,1,8,27,0,0,0,
17,0,7,2,24,1,0,15,3,17,0,2,0,0,
25,19,29,27,26,0,27,0,24,6,15,0,0,0,
7,0,5,19,10,0,25,0,14,10,0,8,0,0,
4,18,10,22,0,6,0,29,28,0,7,22,0,0,
9,15,23,23,5,0,28,18,0,17,0,17,0,0,
19,22,9,5,0,5,0,2,25,16,0,7,0,0,
9,16,23,24,6,0,29,19,0,18,0,18,0,0,
25,5,9,19,17,0,0,15,25,1,0,8,0,0,
17,29,21,24,16,0,16,12,0,27,19,0,0,0,
20,28,0,7,5,0,19,0,16,5,1,0,0,0,
2,5,3,0,14,15,0,2,25,9,0,11,0,0,
12,12,26,0,13,9,20,0,26,0,21,6,0,0,
18,9,10,17,23,0,18,22,0,25,3,0,0,0,
16,1,2,15,26,0,5,17,0,0,3,0,0,0,
25,27,26,16,21,0,8,4,0,14,2,0,0,0,
27,0,23,11,3,22,0,27,16,16,0,18,0,0,
9,3,26,2,0,3,0,2,16,26,0,13,0,0,
2,5,3,0,14,16,0,2,25,9,0,11,0,0,
18,8,0,2,24,1,0,16,3,17,0,3,0,0,
9,3,26,1,0,2,0,1,15,25,0,13,0,0,
25,19,0,27,26,0,27,0,24,6,16,0,0,0,
15,7,18,24,16,0,17,23,0,0,9,1,0,0,
0,23,29,26,3,15,0,7,12,0,2,15,0,0,
27,24,0,11,3,22,0,27,16,16,0,18,0,0,
0,5,18,13,14,22,0,15,26,0,16,7,0,0,
4,0,17,2,15,27,28,7,0,0,29,15,0,0,
25,5,9,19,16,0,0,14,25,1,0,8,0,0,
		others => 0);
	end function;
end package body;
