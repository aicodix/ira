-- code table generated from table_scalar.txt by generate_table_scalar_vhd.cc
--
-- Copyright 2019 Ahmet Inan <inan@aicodix.de>

use work.ldpc_scalar.all;

package table_scalar is
	function init_scalar_parities return scalar_parities;
	function init_scalar_counts return scalar_counts;
	function init_scalar_offsets return scalar_offsets;
end package;

package body table_scalar is
	function init_scalar_parities return scalar_parities is
	begin
		return 2880;
	end function;

	function init_scalar_counts return scalar_counts is
	begin
		return (
15,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
16,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
18,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
19,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
17,
		others => count_scalar'low);
	end function;

	function init_scalar_offsets return scalar_offsets is
	begin
		return (
77,927,1800,1896,3082,4680,5548,5622,7560,7888,9430,10440,12301,13107,13320,
78,928,1801,1897,3083,4681,5549,5623,7561,7889,9431,10441,12302,13108,13321,15840,
79,929,1802,1898,3084,4682,5550,5624,7562,7890,9432,10442,12303,13109,13322,15841,
80,930,1803,1899,3085,4683,5551,5625,7563,7891,9433,10443,12304,13110,13323,15842,
81,931,1804,1900,3086,4684,5552,5626,7564,7892,9434,10444,12305,13111,13324,15843,
82,932,1805,1901,3087,4685,5553,5627,7565,7893,9435,10445,12306,13112,13325,15844,
83,933,1806,1902,3088,4686,5554,5628,7566,7894,9436,10446,12307,13113,13326,15845,
84,934,1807,1903,3089,4687,5555,5629,7567,7895,9437,10447,12308,13114,13327,15846,
85,935,1808,1904,3090,4688,5556,5630,7568,7896,9438,10448,12309,13115,13328,15847,
86,936,1809,1905,3091,4689,5557,5631,7569,7897,9439,10449,12310,13116,13329,15848,
87,937,1810,1906,3092,4690,5558,5632,7570,7898,9440,10450,12311,13117,13330,15849,
88,938,1811,1907,3093,4691,5559,5633,7571,7899,9441,10451,12312,13118,13331,15850,
89,939,1812,1908,3094,4692,5560,5634,7572,7900,9442,10452,12313,13119,13332,15851,
90,940,1813,1909,3095,4693,5561,5635,7573,7901,9443,10453,12314,13120,13333,15852,
91,941,1814,1910,3096,4694,5562,5636,7574,7902,9444,10454,12315,13121,13334,15853,
92,942,1815,1911,3097,4695,5563,5637,7575,7903,9445,10455,12316,13122,13335,15854,
93,943,1816,1912,3098,4696,5564,5638,7576,7904,9446,10456,12317,13123,13336,15855,
94,944,1817,1913,3099,4697,5565,5639,7577,7905,9447,10457,12318,13124,13337,15856,
95,945,1818,1914,3100,4698,5566,5640,7578,7906,9448,10458,12319,13125,13338,15857,
96,946,1819,1915,3101,4699,5567,5641,7579,7907,9449,10459,12320,13126,13339,15858,
97,947,1820,1916,3102,4700,5568,5642,7580,7908,9450,10460,12321,13127,13340,15859,
98,948,1821,1917,3103,4701,5569,5643,7581,7909,9451,10461,12322,13128,13341,15860,
99,949,1822,1918,3104,4702,5570,5644,7582,7910,9452,10462,12323,13129,13342,15861,
100,950,1823,1919,3105,4703,5571,5645,7583,7911,9453,10463,12324,13130,13343,15862,
101,951,1824,1920,3106,4704,5572,5646,7584,7912,9454,10464,12325,13131,13344,15863,
102,952,1825,1921,3107,4705,5573,5647,7585,7913,9455,10465,12326,13132,13345,15864,
103,953,1826,1922,3108,4706,5574,5648,7586,7914,9456,10466,12327,13133,13346,15865,
104,954,1827,1923,3109,4707,5575,5649,7587,7915,9457,10467,12328,13134,13347,15866,
105,955,1828,1924,3110,4708,5576,5650,7588,7916,9458,10468,12329,13135,13348,15867,
106,956,1829,1925,3111,4709,5577,5651,7589,7917,9459,10469,12330,13136,13349,15868,
107,957,1830,1926,3112,4710,5578,5652,7590,7918,9460,10470,12331,13137,13350,15869,
108,958,1831,1927,3113,4711,5579,5653,7591,7919,9461,10471,12332,13138,13351,15870,
109,959,1832,1928,3114,4712,5580,5654,7560,7592,9462,10472,12333,13139,13352,15871,
110,960,1833,1929,3115,4713,5581,5655,7561,7593,9463,10473,12334,13140,13353,15872,
111,961,1834,1930,3116,4714,5582,5656,7562,7594,9464,10474,12335,13141,13354,15873,
112,962,1835,1931,3117,4715,5583,5657,7563,7595,9465,10475,12336,13142,13355,15874,
113,963,1836,1932,3118,4716,5584,5658,7564,7596,9466,10476,12337,13143,13356,15875,
114,964,1837,1933,3119,4717,5585,5659,7565,7597,9467,10477,12338,13144,13357,15876,
115,965,1838,1934,3120,4718,5586,5660,7566,7598,9468,10478,12339,13145,13358,15877,
116,966,1839,1935,3121,4719,5587,5661,7567,7599,9469,10479,12340,13146,13359,15878,
117,967,1840,1936,3122,4720,5588,5662,7568,7600,9470,10480,12341,13147,13360,15879,
118,968,1841,1937,3123,4721,5589,5663,7569,7601,9471,10481,12342,13148,13361,15880,
119,969,1842,1938,3124,4722,5590,5664,7570,7602,9472,10482,12343,13149,13362,15881,
120,970,1843,1939,3125,4723,5591,5665,7571,7603,9473,10483,12344,13150,13363,15882,
121,971,1844,1940,3126,4724,5592,5666,7572,7604,9474,10484,12345,13151,13364,15883,
122,972,1845,1941,3127,4725,5593,5667,7573,7605,9475,10485,12346,13152,13365,15884,
123,973,1846,1942,3128,4726,5594,5668,7574,7606,9476,10486,12347,13153,13366,15885,
124,974,1847,1943,3129,4727,5595,5669,7575,7607,9477,10487,12348,13154,13367,15886,
125,975,1848,1944,3130,4728,5596,5670,7576,7608,9478,10488,12349,13155,13368,15887,
126,976,1849,1945,3131,4729,5597,5671,7577,7609,9479,10489,12350,13156,13369,15888,
127,977,1850,1946,3132,4730,5598,5672,7578,7610,9480,10490,12351,13157,13370,15889,
128,978,1851,1947,3133,4731,5599,5673,7579,7611,9481,10491,12352,13158,13371,15890,
129,979,1852,1948,3134,4732,5600,5674,7580,7612,9482,10492,12353,13159,13372,15891,
130,980,1853,1949,3135,4733,5601,5675,7581,7613,9483,10493,12354,13160,13373,15892,
131,981,1854,1950,3136,4734,5602,5676,7582,7614,9484,10494,12355,13161,13374,15893,
132,982,1855,1951,3137,4735,5603,5677,7583,7615,9485,10495,12356,13162,13375,15894,
133,983,1856,1952,3138,4736,5604,5678,7584,7616,9486,10496,12357,13163,13376,15895,
134,984,1857,1953,3139,4737,5605,5679,7585,7617,9487,10497,12358,13164,13377,15896,
135,985,1858,1954,3140,4738,5606,5680,7586,7618,9488,10498,12359,13165,13378,15897,
136,986,1859,1955,3141,4739,5607,5681,7587,7619,9489,10499,12360,13166,13379,15898,
137,987,1860,1956,3142,4740,5608,5682,7588,7620,9490,10500,12361,13167,13380,15899,
138,988,1861,1957,3143,4741,5609,5683,7589,7621,9491,10501,12362,13168,13381,15900,
139,989,1862,1958,3144,4742,5610,5684,7590,7622,9492,10502,12363,13169,13382,15901,
140,990,1863,1959,3145,4743,5611,5685,7591,7623,9493,10503,12364,13170,13383,15902,
141,991,1864,1960,3146,4744,5612,5686,7592,7624,9494,10504,12365,13171,13384,15903,
142,992,1865,1961,3147,4745,5613,5687,7593,7625,9495,10505,12366,13172,13385,15904,
143,993,1866,1962,3148,4746,5614,5688,7594,7626,9496,10506,12367,13173,13386,15905,
144,994,1867,1963,3149,4747,5615,5689,7595,7627,9497,10507,12368,13174,13387,15906,
145,995,1868,1964,3150,4748,5616,5690,7596,7628,9498,10508,12369,13175,13388,15907,
146,996,1869,1965,3151,4749,5617,5691,7597,7629,9499,10509,12370,13176,13389,15908,
147,997,1870,1966,3152,4750,5618,5692,7598,7630,9500,10510,12371,13177,13390,15909,
148,998,1871,1967,3153,4751,5619,5693,7599,7631,9501,10511,12372,13178,13391,15910,
149,999,1872,1968,3154,4752,5620,5694,7600,7632,9502,10512,12373,13179,13392,15911,
150,1000,1873,1969,3155,4753,5621,5695,7601,7633,9503,10513,12374,13180,13393,15912,
151,1001,1874,1970,3156,4754,5622,5696,7602,7634,9504,10514,12375,13181,13394,15913,
152,1002,1875,1971,3157,4755,5623,5697,7603,7635,9505,10515,12376,13182,13395,15914,
153,1003,1876,1972,3158,4756,5624,5698,7604,7636,9506,10516,12377,13183,13396,15915,
154,1004,1877,1973,3159,4757,5625,5699,7605,7637,9507,10517,12378,13184,13397,15916,
155,1005,1878,1974,3160,4758,5626,5700,7606,7638,9508,10518,12379,13185,13398,15917,
156,1006,1879,1975,3161,4759,5627,5701,7607,7639,9509,10519,12380,13186,13399,15918,
157,1007,1880,1976,3162,4760,5628,5702,7608,7640,9510,10520,12381,13187,13400,15919,
158,1008,1881,1977,3163,4761,5629,5703,7609,7641,9511,10521,12382,13188,13401,15920,
159,1009,1882,1978,3164,4762,5630,5704,7610,7642,9512,10522,12383,13189,13402,15921,
160,1010,1883,1979,3165,4763,5631,5705,7611,7643,9513,10523,12384,13190,13403,15922,
161,1011,1884,1980,3166,4764,5632,5706,7612,7644,9514,10524,12385,13191,13404,15923,
162,1012,1885,1981,3167,4765,5633,5707,7613,7645,9515,10525,12386,13192,13405,15924,
163,1013,1886,1982,3168,4766,5634,5708,7614,7646,9516,10526,12387,13193,13406,15925,
164,1014,1887,1983,3169,4767,5635,5709,7615,7647,9517,10527,12388,13194,13407,15926,
165,1015,1888,1984,3170,4768,5636,5710,7616,7648,9518,10528,12389,13195,13408,15927,
166,1016,1889,1985,3171,4769,5637,5711,7617,7649,9519,10529,12390,13196,13409,15928,
167,1017,1890,1986,3172,4770,5638,5712,7618,7650,9520,10530,12391,13197,13410,15929,
168,1018,1891,1987,3173,4771,5639,5713,7619,7651,9521,10531,12392,13198,13411,15930,
169,1019,1892,1988,3174,4772,5640,5714,7620,7652,9522,10532,12393,13199,13412,15931,
170,1020,1893,1989,3175,4773,5641,5715,7621,7653,9523,10533,12394,13200,13413,15932,
171,1021,1894,1990,3176,4774,5642,5716,7622,7654,9524,10534,12395,13201,13414,15933,
172,1022,1895,1991,3177,4775,5643,5717,7623,7655,9525,10535,12396,13202,13415,15934,
173,1023,1896,1992,3178,4776,5644,5718,7624,7656,9526,10536,12397,13203,13416,15935,
174,1024,1897,1993,3179,4777,5645,5719,7625,7657,9527,10537,12398,13204,13417,15936,
175,1025,1898,1994,3180,4778,5646,5720,7626,7658,9528,10538,12399,13205,13418,15937,
176,1026,1899,1995,3181,4779,5647,5721,7627,7659,9529,10539,12400,13206,13419,15938,
177,1027,1900,1996,3182,4780,5648,5722,7628,7660,9530,10540,12401,13207,13420,15939,
178,1028,1901,1997,3183,4781,5649,5723,7629,7661,9531,10541,12402,13208,13421,15940,
179,1029,1902,1998,3184,4782,5650,5724,7630,7662,9532,10542,12403,13209,13422,15941,
180,1030,1903,1999,3185,4783,5651,5725,7631,7663,9533,10543,12404,13210,13423,15942,
181,1031,1904,2000,3186,4784,5652,5726,7632,7664,9534,10544,12405,13211,13424,15943,
182,1032,1905,2001,3187,4785,5653,5727,7633,7665,9535,10545,12406,13212,13425,15944,
183,1033,1906,2002,3188,4786,5654,5728,7634,7666,9536,10546,12407,13213,13426,15945,
184,1034,1907,2003,3189,4787,5655,5729,7635,7667,9537,10547,12408,13214,13427,15946,
185,1035,1908,2004,3190,4788,5656,5730,7636,7668,9538,10548,12409,13215,13428,15947,
186,1036,1909,2005,3191,4789,5657,5731,7637,7669,9539,10549,12410,13216,13429,15948,
187,1037,1910,2006,3192,4790,5658,5732,7638,7670,9540,10550,12411,13217,13430,15949,
188,1038,1911,2007,3193,4791,5659,5733,7639,7671,9541,10551,12412,13218,13431,15950,
189,1039,1912,2008,3194,4792,5660,5734,7640,7672,9542,10552,12413,13219,13432,15951,
190,1040,1913,2009,3195,4793,5661,5735,7641,7673,9543,10553,12414,13220,13433,15952,
191,1041,1914,2010,3196,4794,5662,5736,7642,7674,9544,10554,12415,13221,13434,15953,
192,1042,1915,2011,3197,4795,5663,5737,7643,7675,9545,10555,12416,13222,13435,15954,
193,1043,1916,2012,3198,4796,5664,5738,7644,7676,9546,10556,12417,13223,13436,15955,
194,1044,1917,2013,3199,4797,5665,5739,7645,7677,9547,10557,12418,13224,13437,15956,
195,1045,1918,2014,3200,4798,5666,5740,7646,7678,9548,10558,12419,13225,13438,15957,
196,1046,1919,2015,3201,4799,5667,5741,7647,7679,9549,10559,12420,13226,13439,15958,
197,1047,1920,2016,3202,4800,5668,5742,7648,7680,9550,10560,12421,13227,13440,15959,
198,1048,1921,2017,3203,4801,5669,5743,7649,7681,9551,10561,12422,13228,13441,15960,
199,1049,1922,2018,3204,4802,5670,5744,7650,7682,9552,10562,12423,13229,13442,15961,
200,1050,1923,2019,3205,4803,5671,5745,7651,7683,9553,10563,12424,13230,13443,15962,
201,1051,1924,2020,3206,4804,5672,5746,7652,7684,9554,10564,12425,13231,13444,15963,
202,1052,1925,2021,3207,4805,5673,5747,7653,7685,9555,10565,12426,13232,13445,15964,
203,1053,1926,2022,3208,4806,5674,5748,7654,7686,9556,10566,12427,13233,13446,15965,
204,1054,1927,2023,3209,4807,5675,5749,7655,7687,9557,10567,12428,13234,13447,15966,
205,1055,1928,2024,3210,4808,5676,5750,7656,7688,9558,10568,12429,13235,13448,15967,
206,1056,1929,2025,3211,4809,5677,5751,7657,7689,9559,10569,12430,13236,13449,15968,
207,1057,1930,2026,3212,4810,5678,5752,7658,7690,9560,10570,12431,13237,13450,15969,
208,1058,1931,2027,3213,4811,5679,5753,7659,7691,9561,10571,12432,13238,13451,15970,
209,1059,1932,2028,3214,4812,5680,5754,7660,7692,9562,10572,12433,13239,13452,15971,
210,1060,1933,2029,3215,4813,5681,5755,7661,7693,9563,10573,12434,13240,13453,15972,
211,1061,1934,2030,3216,4814,5682,5756,7662,7694,9564,10574,12435,13241,13454,15973,
212,1062,1935,2031,3217,4815,5683,5757,7663,7695,9565,10575,12436,13242,13455,15974,
213,1063,1936,2032,3218,4816,5684,5758,7664,7696,9566,10576,12437,13243,13456,15975,
214,1064,1937,2033,3219,4817,5685,5759,7665,7697,9567,10577,12438,13244,13457,15976,
215,1065,1938,2034,3220,4818,5400,5686,7666,7698,9568,10578,12439,13245,13458,15977,
216,1066,1939,2035,3221,4819,5401,5687,7667,7699,9569,10579,12440,13246,13459,15978,
217,1067,1940,2036,3222,4820,5402,5688,7668,7700,9570,10580,12441,13247,13460,15979,
218,1068,1941,2037,3223,4821,5403,5689,7669,7701,9571,10581,12442,13248,13461,15980,
219,1069,1942,2038,3224,4822,5404,5690,7670,7702,9572,10582,12443,13249,13462,15981,
220,1070,1943,2039,3225,4823,5405,5691,7671,7703,9573,10583,12444,13250,13463,15982,
221,1071,1944,2040,3226,4824,5406,5692,7672,7704,9574,10584,12445,13251,13464,15983,
222,1072,1945,2041,3227,4825,5407,5693,7673,7705,9575,10585,12446,13252,13465,15984,
223,1073,1946,2042,3228,4826,5408,5694,7674,7706,9576,10586,12447,13253,13466,15985,
224,1074,1947,2043,3229,4827,5409,5695,7675,7707,9577,10587,12448,13254,13467,15986,
225,1075,1948,2044,3230,4828,5410,5696,7676,7708,9578,10588,12449,13255,13468,15987,
226,1076,1949,2045,3231,4829,5411,5697,7677,7709,9579,10589,12450,13256,13469,15988,
227,1077,1950,2046,3232,4830,5412,5698,7678,7710,9580,10590,12451,13257,13470,15989,
228,1078,1951,2047,3233,4831,5413,5699,7679,7711,9581,10591,12452,13258,13471,15990,
229,1079,1952,2048,3234,4832,5414,5700,7680,7712,9582,10592,12453,13259,13472,15991,
230,720,1953,2049,3235,4833,5415,5701,7681,7713,9583,10593,12454,13260,13473,15992,
231,721,1954,2050,3236,4834,5416,5702,7682,7714,9584,10594,12455,13261,13474,15993,
232,722,1955,2051,3237,4835,5417,5703,7683,7715,9585,10595,12456,13262,13475,15994,
233,723,1956,2052,3238,4836,5418,5704,7684,7716,9586,10596,12457,13263,13476,15995,
234,724,1957,2053,3239,4837,5419,5705,7685,7717,9587,10597,12458,13264,13477,15996,
235,725,1958,2054,2880,4838,5420,5706,7686,7718,9588,10598,12459,13265,13478,15997,
236,726,1959,2055,2881,4839,5421,5707,7687,7719,9589,10599,12460,13266,13479,15998,
237,727,1960,2056,2882,4840,5422,5708,7688,7720,9590,10600,12461,13267,13480,15999,
238,728,1961,2057,2883,4841,5423,5709,7689,7721,9591,10601,12462,13268,13481,16000,
239,729,1962,2058,2884,4842,5424,5710,7690,7722,9592,10602,12463,13269,13482,16001,
240,730,1963,2059,2885,4843,5425,5711,7691,7723,9593,10603,12464,13270,13483,16002,
241,731,1964,2060,2886,4844,5426,5712,7692,7724,9594,10604,12465,13271,13484,16003,
242,732,1965,2061,2887,4845,5427,5713,7693,7725,9595,10605,12466,13272,13485,16004,
243,733,1966,2062,2888,4846,5428,5714,7694,7726,9596,10606,12467,13273,13486,16005,
244,734,1967,2063,2889,4847,5429,5715,7695,7727,9597,10607,12468,13274,13487,16006,
245,735,1968,2064,2890,4848,5430,5716,7696,7728,9598,10608,12469,13275,13488,16007,
246,736,1969,2065,2891,4849,5431,5717,7697,7729,9599,10609,12470,13276,13489,16008,
247,737,1970,2066,2892,4850,5432,5718,7698,7730,9600,10610,12471,13277,13490,16009,
248,738,1971,2067,2893,4851,5433,5719,7699,7731,9601,10611,12472,13278,13491,16010,
249,739,1972,2068,2894,4852,5434,5720,7700,7732,9602,10612,12473,13279,13492,16011,
250,740,1973,2069,2895,4853,5435,5721,7701,7733,9603,10613,12474,13280,13493,16012,
251,741,1974,2070,2896,4854,5436,5722,7702,7734,9604,10614,12475,13281,13494,16013,
252,742,1975,2071,2897,4855,5437,5723,7703,7735,9605,10615,12476,13282,13495,16014,
253,743,1976,2072,2898,4856,5438,5724,7704,7736,9606,10616,12477,13283,13496,16015,
254,744,1977,2073,2899,4857,5439,5725,7705,7737,9607,10617,12478,13284,13497,16016,
255,745,1978,2074,2900,4858,5440,5726,7706,7738,9608,10618,12479,13285,13498,16017,
256,746,1979,2075,2901,4859,5441,5727,7707,7739,9609,10619,12480,13286,13499,16018,
257,747,1980,2076,2902,4860,5442,5728,7708,7740,9610,10620,12481,13287,13500,16019,
258,748,1981,2077,2903,4861,5443,5729,7709,7741,9611,10621,12482,13288,13501,16020,
259,749,1982,2078,2904,4862,5444,5730,7710,7742,9612,10622,12483,13289,13502,16021,
260,750,1983,2079,2905,4863,5445,5731,7711,7743,9613,10623,12484,13290,13503,16022,
261,751,1984,2080,2906,4864,5446,5732,7712,7744,9614,10624,12485,13291,13504,16023,
262,752,1985,2081,2907,4865,5447,5733,7713,7745,9615,10625,12486,13292,13505,16024,
263,753,1986,2082,2908,4866,5448,5734,7714,7746,9616,10626,12487,13293,13506,16025,
264,754,1987,2083,2909,4867,5449,5735,7715,7747,9617,10627,12488,13294,13507,16026,
265,755,1988,2084,2910,4868,5450,5736,7716,7748,9618,10628,12489,13295,13508,16027,
266,756,1989,2085,2911,4869,5451,5737,7717,7749,9619,10629,12490,13296,13509,16028,
267,757,1990,2086,2912,4870,5452,5738,7718,7750,9620,10630,12491,13297,13510,16029,
268,758,1991,2087,2913,4871,5453,5739,7719,7751,9621,10631,12492,13298,13511,16030,
269,759,1992,2088,2914,4872,5454,5740,7720,7752,9622,10632,12493,13299,13512,16031,
270,760,1993,2089,2915,4873,5455,5741,7721,7753,9623,10633,12494,13300,13513,16032,
271,761,1994,2090,2916,4874,5456,5742,7722,7754,9624,10634,12495,13301,13514,16033,
272,762,1995,2091,2917,4875,5457,5743,7723,7755,9625,10635,12496,13302,13515,16034,
273,763,1996,2092,2918,4876,5458,5744,7724,7756,9626,10636,12497,13303,13516,16035,
274,764,1997,2093,2919,4877,5459,5745,7725,7757,9627,10637,12498,13304,13517,16036,
275,765,1998,2094,2920,4878,5460,5746,7726,7758,9628,10638,12499,13305,13518,16037,
276,766,1999,2095,2921,4879,5461,5747,7727,7759,9629,10639,12500,13306,13519,16038,
277,767,2000,2096,2922,4880,5462,5748,7728,7760,9630,10640,12501,13307,13520,16039,
278,768,2001,2097,2923,4881,5463,5749,7729,7761,9631,10641,12502,13308,13521,16040,
279,769,2002,2098,2924,4882,5464,5750,7730,7762,9632,10642,12503,13309,13522,16041,
280,770,2003,2099,2925,4883,5465,5751,7731,7763,9633,10643,12504,13310,13523,16042,
281,771,2004,2100,2926,4884,5466,5752,7732,7764,9634,10644,12505,13311,13524,16043,
282,772,2005,2101,2927,4885,5467,5753,7733,7765,9635,10645,12506,13312,13525,16044,
283,773,2006,2102,2928,4886,5468,5754,7734,7766,9636,10646,12507,13313,13526,16045,
284,774,2007,2103,2929,4887,5469,5755,7735,7767,9637,10647,12508,13314,13527,16046,
285,775,2008,2104,2930,4888,5470,5756,7736,7768,9638,10648,12509,13315,13528,16047,
286,776,2009,2105,2931,4889,5471,5757,7737,7769,9639,10649,12510,13316,13529,16048,
287,777,2010,2106,2932,4890,5472,5758,7738,7770,9640,10650,12511,13317,13530,16049,
288,778,2011,2107,2933,4891,5473,5759,7739,7771,9641,10651,12512,13318,13531,16050,
289,779,2012,2108,2934,4892,5400,5474,7740,7772,9642,10652,12513,13319,13532,16051,
290,780,2013,2109,2935,4893,5401,5475,7741,7773,9643,10653,12514,12960,13533,16052,
291,781,2014,2110,2936,4894,5402,5476,7742,7774,9644,10654,12515,12961,13534,16053,
292,782,2015,2111,2937,4895,5403,5477,7743,7775,9645,10655,12516,12962,13535,16054,
293,783,2016,2112,2938,4896,5404,5478,7744,7776,9646,10656,12517,12963,13536,16055,
294,784,2017,2113,2939,4897,5405,5479,7745,7777,9647,10657,12518,12964,13537,16056,
295,785,2018,2114,2940,4898,5406,5480,7746,7778,9648,10658,12519,12965,13538,16057,
296,786,2019,2115,2941,4899,5407,5481,7747,7779,9649,10659,12520,12966,13539,16058,
297,787,2020,2116,2942,4900,5408,5482,7748,7780,9650,10660,12521,12967,13540,16059,
298,788,2021,2117,2943,4901,5409,5483,7749,7781,9651,10661,12522,12968,13541,16060,
299,789,2022,2118,2944,4902,5410,5484,7750,7782,9652,10662,12523,12969,13542,16061,
300,790,2023,2119,2945,4903,5411,5485,7751,7783,9653,10663,12524,12970,13543,16062,
301,791,2024,2120,2946,4904,5412,5486,7752,7784,9654,10664,12525,12971,13544,16063,
302,792,2025,2121,2947,4905,5413,5487,7753,7785,9655,10665,12526,12972,13545,16064,
303,793,2026,2122,2948,4906,5414,5488,7754,7786,9656,10666,12527,12973,13546,16065,
304,794,2027,2123,2949,4907,5415,5489,7755,7787,9657,10667,12528,12974,13547,16066,
305,795,2028,2124,2950,4908,5416,5490,7756,7788,9658,10668,12529,12975,13548,16067,
306,796,2029,2125,2951,4909,5417,5491,7757,7789,9659,10669,12530,12976,13549,16068,
307,797,2030,2126,2952,4910,5418,5492,7758,7790,9660,10670,12531,12977,13550,16069,
308,798,2031,2127,2953,4911,5419,5493,7759,7791,9661,10671,12532,12978,13551,16070,
309,799,2032,2128,2954,4912,5420,5494,7760,7792,9662,10672,12533,12979,13552,16071,
310,800,2033,2129,2955,4913,5421,5495,7761,7793,9663,10673,12534,12980,13553,16072,
311,801,2034,2130,2956,4914,5422,5496,7762,7794,9664,10674,12535,12981,13554,16073,
312,802,2035,2131,2957,4915,5423,5497,7763,7795,9665,10675,12536,12982,13555,16074,
313,803,2036,2132,2958,4916,5424,5498,7764,7796,9666,10676,12537,12983,13556,16075,
314,804,2037,2133,2959,4917,5425,5499,7765,7797,9667,10677,12538,12984,13557,16076,
315,805,2038,2134,2960,4918,5426,5500,7766,7798,9668,10678,12539,12985,13558,16077,
316,806,2039,2135,2961,4919,5427,5501,7767,7799,9669,10679,12540,12986,13559,16078,
317,807,2040,2136,2962,4920,5428,5502,7768,7800,9670,10680,12541,12987,13560,16079,
318,808,2041,2137,2963,4921,5429,5503,7769,7801,9671,10681,12542,12988,13561,16080,
319,809,2042,2138,2964,4922,5430,5504,7770,7802,9672,10682,12543,12989,13562,16081,
320,810,2043,2139,2965,4923,5431,5505,7771,7803,9673,10683,12544,12990,13563,16082,
321,811,2044,2140,2966,4924,5432,5506,7772,7804,9674,10684,12545,12991,13564,16083,
322,812,2045,2141,2967,4925,5433,5507,7773,7805,9675,10685,12546,12992,13565,16084,
323,813,2046,2142,2968,4926,5434,5508,7774,7806,9676,10686,12547,12993,13566,16085,
324,814,2047,2143,2969,4927,5435,5509,7775,7807,9677,10687,12548,12994,13567,16086,
325,815,2048,2144,2970,4928,5436,5510,7776,7808,9678,10688,12549,12995,13568,16087,
326,816,2049,2145,2971,4929,5437,5511,7777,7809,9679,10689,12550,12996,13569,16088,
327,817,2050,2146,2972,4930,5438,5512,7778,7810,9680,10690,12551,12997,13570,16089,
328,818,2051,2147,2973,4931,5439,5513,7779,7811,9681,10691,12552,12998,13571,16090,
329,819,2052,2148,2974,4932,5440,5514,7780,7812,9682,10692,12553,12999,13572,16091,
330,820,2053,2149,2975,4933,5441,5515,7781,7813,9683,10693,12554,13000,13573,16092,
331,821,2054,2150,2976,4934,5442,5516,7782,7814,9684,10694,12555,13001,13574,16093,
332,822,2055,2151,2977,4935,5443,5517,7783,7815,9685,10695,12556,13002,13575,16094,
333,823,2056,2152,2978,4936,5444,5518,7784,7816,9686,10696,12557,13003,13576,16095,
334,824,2057,2153,2979,4937,5445,5519,7785,7817,9687,10697,12558,13004,13577,16096,
335,825,2058,2154,2980,4938,5446,5520,7786,7818,9688,10698,12559,13005,13578,16097,
336,826,2059,2155,2981,4939,5447,5521,7787,7819,9689,10699,12560,13006,13579,16098,
337,827,2060,2156,2982,4940,5448,5522,7788,7820,9690,10700,12561,13007,13580,16099,
338,828,2061,2157,2983,4941,5449,5523,7789,7821,9691,10701,12562,13008,13581,16100,
339,829,2062,2158,2984,4942,5450,5524,7790,7822,9692,10702,12563,13009,13582,16101,
340,830,2063,2159,2985,4943,5451,5525,7791,7823,9693,10703,12564,13010,13583,16102,
341,831,1800,2064,2986,4944,5452,5526,7792,7824,9694,10704,12565,13011,13584,16103,
342,832,1801,2065,2987,4945,5453,5527,7793,7825,9695,10705,12566,13012,13585,16104,
343,833,1802,2066,2988,4946,5454,5528,7794,7826,9696,10706,12567,13013,13586,16105,
344,834,1803,2067,2989,4947,5455,5529,7795,7827,9697,10707,12568,13014,13587,16106,
345,835,1804,2068,2990,4948,5456,5530,7796,7828,9698,10708,12569,13015,13588,16107,
346,836,1805,2069,2991,4949,5457,5531,7797,7829,9699,10709,12570,13016,13589,16108,
347,837,1806,2070,2992,4950,5458,5532,7798,7830,9700,10710,12571,13017,13590,16109,
348,838,1807,2071,2993,4951,5459,5533,7799,7831,9701,10711,12572,13018,13591,16110,
349,839,1808,2072,2994,4952,5460,5534,7800,7832,9702,10712,12573,13019,13592,16111,
350,840,1809,2073,2995,4953,5461,5535,7801,7833,9703,10713,12574,13020,13593,16112,
351,841,1810,2074,2996,4954,5462,5536,7802,7834,9704,10714,12575,13021,13594,16113,
352,842,1811,2075,2997,4955,5463,5537,7803,7835,9705,10715,12576,13022,13595,16114,
353,843,1812,2076,2998,4956,5464,5538,7804,7836,9706,10716,12577,13023,13596,16115,
354,844,1813,2077,2999,4957,5465,5539,7805,7837,9707,10717,12578,13024,13597,16116,
355,845,1814,2078,3000,4958,5466,5540,7806,7838,9708,10718,12579,13025,13598,16117,
356,846,1815,2079,3001,4959,5467,5541,7807,7839,9709,10719,12580,13026,13599,16118,
357,847,1816,2080,3002,4960,5468,5542,7808,7840,9710,10720,12581,13027,13600,16119,
358,848,1817,2081,3003,4961,5469,5543,7809,7841,9711,10721,12582,13028,13601,16120,
359,849,1818,2082,3004,4962,5470,5544,7810,7842,9712,10722,12583,13029,13602,16121,
0,850,1819,2083,3005,4963,5471,5545,7811,7843,9713,10723,12584,13030,13603,16122,
1,851,1820,2084,3006,4964,5472,5546,7812,7844,9714,10724,12585,13031,13604,16123,
2,852,1821,2085,3007,4965,5473,5547,7813,7845,9715,10725,12586,13032,13605,16124,
3,853,1822,2086,3008,4966,5474,5548,7814,7846,9716,10726,12587,13033,13606,16125,
4,854,1823,2087,3009,4967,5475,5549,7815,7847,9717,10727,12588,13034,13607,16126,
5,855,1824,2088,3010,4968,5476,5550,7816,7848,9718,10728,12589,13035,13608,16127,
6,856,1825,2089,3011,4969,5477,5551,7817,7849,9719,10729,12590,13036,13609,16128,
7,857,1826,2090,3012,4970,5478,5552,7818,7850,9360,10730,12591,13037,13610,16129,
8,858,1827,2091,3013,4971,5479,5553,7819,7851,9361,10731,12592,13038,13611,16130,
9,859,1828,2092,3014,4972,5480,5554,7820,7852,9362,10732,12593,13039,13612,16131,
10,860,1829,2093,3015,4973,5481,5555,7821,7853,9363,10733,12594,13040,13613,16132,
11,861,1830,2094,3016,4974,5482,5556,7822,7854,9364,10734,12595,13041,13614,16133,
12,862,1831,2095,3017,4975,5483,5557,7823,7855,9365,10735,12596,13042,13615,16134,
13,863,1832,2096,3018,4976,5484,5558,7824,7856,9366,10736,12597,13043,13616,16135,
14,864,1833,2097,3019,4977,5485,5559,7825,7857,9367,10737,12598,13044,13617,16136,
15,865,1834,2098,3020,4978,5486,5560,7826,7858,9368,10738,12599,13045,13618,16137,
16,866,1835,2099,3021,4979,5487,5561,7827,7859,9369,10739,12240,13046,13619,16138,
17,867,1836,2100,3022,4980,5488,5562,7828,7860,9370,10740,12241,13047,13620,16139,
18,868,1837,2101,3023,4981,5489,5563,7829,7861,9371,10741,12242,13048,13621,16140,
19,869,1838,2102,3024,4982,5490,5564,7830,7862,9372,10742,12243,13049,13622,16141,
20,870,1839,2103,3025,4983,5491,5565,7831,7863,9373,10743,12244,13050,13623,16142,
21,871,1840,2104,3026,4984,5492,5566,7832,7864,9374,10744,12245,13051,13624,16143,
22,872,1841,2105,3027,4985,5493,5567,7833,7865,9375,10745,12246,13052,13625,16144,
23,873,1842,2106,3028,4986,5494,5568,7834,7866,9376,10746,12247,13053,13626,16145,
24,874,1843,2107,3029,4987,5495,5569,7835,7867,9377,10747,12248,13054,13627,16146,
25,875,1844,2108,3030,4988,5496,5570,7836,7868,9378,10748,12249,13055,13628,16147,
26,876,1845,2109,3031,4989,5497,5571,7837,7869,9379,10749,12250,13056,13629,16148,
27,877,1846,2110,3032,4990,5498,5572,7838,7870,9380,10750,12251,13057,13630,16149,
28,878,1847,2111,3033,4991,5499,5573,7839,7871,9381,10751,12252,13058,13631,16150,
29,879,1848,2112,3034,4992,5500,5574,7840,7872,9382,10752,12253,13059,13632,16151,
30,880,1849,2113,3035,4993,5501,5575,7841,7873,9383,10753,12254,13060,13633,16152,
31,881,1850,2114,3036,4994,5502,5576,7842,7874,9384,10754,12255,13061,13634,16153,
32,882,1851,2115,3037,4995,5503,5577,7843,7875,9385,10755,12256,13062,13635,16154,
33,883,1852,2116,3038,4996,5504,5578,7844,7876,9386,10756,12257,13063,13636,16155,
34,884,1853,2117,3039,4997,5505,5579,7845,7877,9387,10757,12258,13064,13637,16156,
35,885,1854,2118,3040,4998,5506,5580,7846,7878,9388,10758,12259,13065,13638,16157,
36,886,1855,2119,3041,4999,5507,5581,7847,7879,9389,10759,12260,13066,13639,16158,
37,887,1856,2120,3042,5000,5508,5582,7848,7880,9390,10760,12261,13067,13640,16159,
38,888,1857,2121,3043,5001,5509,5583,7849,7881,9391,10761,12262,13068,13641,16160,
39,889,1858,2122,3044,5002,5510,5584,7850,7882,9392,10762,12263,13069,13642,16161,
40,890,1859,2123,3045,5003,5511,5585,7851,7883,9393,10763,12264,13070,13643,16162,
41,891,1860,2124,3046,5004,5512,5586,7852,7884,9394,10764,12265,13071,13644,16163,
42,892,1861,2125,3047,5005,5513,5587,7853,7885,9395,10765,12266,13072,13645,16164,
43,893,1862,2126,3048,5006,5514,5588,7854,7886,9396,10766,12267,13073,13646,16165,
44,894,1863,2127,3049,5007,5515,5589,7855,7887,9397,10767,12268,13074,13647,16166,
45,895,1864,2128,3050,5008,5516,5590,7856,7888,9398,10768,12269,13075,13648,16167,
46,896,1865,2129,3051,5009,5517,5591,7857,7889,9399,10769,12270,13076,13649,16168,
47,897,1866,2130,3052,5010,5518,5592,7858,7890,9400,10770,12271,13077,13650,16169,
48,898,1867,2131,3053,5011,5519,5593,7859,7891,9401,10771,12272,13078,13651,16170,
49,899,1868,2132,3054,5012,5520,5594,7860,7892,9402,10772,12273,13079,13652,16171,
50,900,1869,2133,3055,5013,5521,5595,7861,7893,9403,10773,12274,13080,13653,16172,
51,901,1870,2134,3056,5014,5522,5596,7862,7894,9404,10774,12275,13081,13654,16173,
52,902,1871,2135,3057,5015,5523,5597,7863,7895,9405,10775,12276,13082,13655,16174,
53,903,1872,2136,3058,5016,5524,5598,7864,7896,9406,10776,12277,13083,13656,16175,
54,904,1873,2137,3059,5017,5525,5599,7865,7897,9407,10777,12278,13084,13657,16176,
55,905,1874,2138,3060,5018,5526,5600,7866,7898,9408,10778,12279,13085,13658,16177,
56,906,1875,2139,3061,5019,5527,5601,7867,7899,9409,10779,12280,13086,13659,16178,
57,907,1876,2140,3062,5020,5528,5602,7868,7900,9410,10780,12281,13087,13660,16179,
58,908,1877,2141,3063,5021,5529,5603,7869,7901,9411,10781,12282,13088,13661,16180,
59,909,1878,2142,3064,5022,5530,5604,7870,7902,9412,10782,12283,13089,13662,16181,
60,910,1879,2143,3065,5023,5531,5605,7871,7903,9413,10783,12284,13090,13663,16182,
61,911,1880,2144,3066,5024,5532,5606,7872,7904,9414,10784,12285,13091,13664,16183,
62,912,1881,2145,3067,5025,5533,5607,7873,7905,9415,10785,12286,13092,13665,16184,
63,913,1882,2146,3068,5026,5534,5608,7874,7906,9416,10786,12287,13093,13666,16185,
64,914,1883,2147,3069,5027,5535,5609,7875,7907,9417,10787,12288,13094,13667,16186,
65,915,1884,2148,3070,5028,5536,5610,7876,7908,9418,10788,12289,13095,13668,16187,
66,916,1885,2149,3071,5029,5537,5611,7877,7909,9419,10789,12290,13096,13669,16188,
67,917,1886,2150,3072,5030,5538,5612,7878,7910,9420,10790,12291,13097,13670,16189,
68,918,1887,2151,3073,5031,5539,5613,7879,7911,9421,10791,12292,13098,13671,16190,
69,919,1888,2152,3074,5032,5540,5614,7880,7912,9422,10792,12293,13099,13672,16191,
70,920,1889,2153,3075,5033,5541,5615,7881,7913,9423,10793,12294,13100,13673,16192,
71,921,1890,2154,3076,5034,5542,5616,7882,7914,9424,10794,12295,13101,13674,16193,
72,922,1891,2155,3077,5035,5543,5617,7883,7915,9425,10795,12296,13102,13675,16194,
73,923,1892,2156,3078,5036,5544,5618,7884,7916,9426,10796,12297,13103,13676,16195,
74,924,1893,2157,3079,5037,5545,5619,7885,7917,9427,10797,12298,13104,13677,16196,
75,925,1894,2158,3080,5038,5546,5620,7886,7918,9428,10798,12299,13105,13678,16197,
76,926,1895,2159,3081,5039,5547,5621,7887,7919,9429,10799,12300,13106,13679,16198,
59,175,2160,2812,4670,5040,5379,7138,7920,8483,8847,10504,10800,11153,13320,13680,
60,176,2161,2813,4671,5041,5380,7139,7921,8484,8848,10505,10801,11154,13321,13681,
61,177,2162,2814,4672,5042,5381,7140,7922,8485,8849,10506,10802,11155,13322,13682,
62,178,2163,2815,4673,5043,5382,7141,7923,8486,8850,10507,10803,11156,13323,13683,
63,179,2164,2816,4674,5044,5383,7142,7924,8487,8851,10508,10804,11157,13324,13684,
64,180,2165,2817,4675,5045,5384,7143,7925,8488,8852,10509,10805,11158,13325,13685,
65,181,2166,2818,4676,5046,5385,7144,7926,8489,8853,10510,10806,11159,13326,13686,
66,182,2167,2819,4677,5047,5386,7145,7927,8490,8854,10511,10800,10807,13327,13687,
67,183,2168,2820,4678,5048,5387,7146,7928,8491,8855,10512,10801,10808,13328,13688,
68,184,2169,2821,4679,5049,5388,7147,7929,8492,8856,10513,10802,10809,13329,13689,
69,185,2170,2822,4320,5050,5389,7148,7930,8493,8857,10514,10803,10810,13330,13690,
70,186,2171,2823,4321,5051,5390,7149,7931,8494,8858,10515,10804,10811,13331,13691,
71,187,2172,2824,4322,5052,5391,7150,7932,8495,8859,10516,10805,10812,13332,13692,
72,188,2173,2825,4323,5053,5392,7151,7933,8496,8860,10517,10806,10813,13333,13693,
73,189,2174,2826,4324,5054,5393,7152,7934,8497,8861,10518,10807,10814,13334,13694,
74,190,2175,2827,4325,5055,5394,7153,7935,8498,8862,10519,10808,10815,13335,13695,
75,191,2176,2828,4326,5056,5395,7154,7936,8499,8863,10520,10809,10816,13336,13696,
76,192,2177,2829,4327,5057,5396,7155,7937,8500,8864,10521,10810,10817,13337,13697,
77,193,2178,2830,4328,5058,5397,7156,7938,8501,8865,10522,10811,10818,13338,13698,
78,194,2179,2831,4329,5059,5398,7157,7939,8502,8866,10523,10812,10819,13339,13699,
79,195,2180,2832,4330,5060,5399,7158,7940,8503,8867,10524,10813,10820,13340,13700,
80,196,2181,2833,4331,5040,5061,7159,7941,8504,8868,10525,10814,10821,13341,13701,
81,197,2182,2834,4332,5041,5062,7160,7942,8505,8869,10526,10815,10822,13342,13702,
82,198,2183,2835,4333,5042,5063,7161,7943,8506,8870,10527,10816,10823,13343,13703,
83,199,2184,2836,4334,5043,5064,7162,7944,8507,8871,10528,10817,10824,13344,13704,
84,200,2185,2837,4335,5044,5065,7163,7945,8508,8872,10529,10818,10825,13345,13705,
85,201,2186,2838,4336,5045,5066,7164,7946,8509,8873,10530,10819,10826,13346,13706,
86,202,2187,2839,4337,5046,5067,7165,7947,8510,8874,10531,10820,10827,13347,13707,
87,203,2188,2840,4338,5047,5068,7166,7948,8511,8875,10532,10821,10828,13348,13708,
88,204,2189,2841,4339,5048,5069,7167,7949,8512,8876,10533,10822,10829,13349,13709,
89,205,2190,2842,4340,5049,5070,7168,7950,8513,8877,10534,10823,10830,13350,13710,
90,206,2191,2843,4341,5050,5071,7169,7951,8514,8878,10535,10824,10831,13351,13711,
91,207,2192,2844,4342,5051,5072,7170,7952,8515,8879,10536,10825,10832,13352,13712,
92,208,2193,2845,4343,5052,5073,7171,7953,8516,8880,10537,10826,10833,13353,13713,
93,209,2194,2846,4344,5053,5074,7172,7954,8517,8881,10538,10827,10834,13354,13714,
94,210,2195,2847,4345,5054,5075,7173,7955,8518,8882,10539,10828,10835,13355,13715,
95,211,2196,2848,4346,5055,5076,7174,7956,8519,8883,10540,10829,10836,13356,13716,
96,212,2197,2849,4347,5056,5077,7175,7957,8520,8884,10541,10830,10837,13357,13717,
97,213,2198,2850,4348,5057,5078,7176,7958,8521,8885,10542,10831,10838,13358,13718,
98,214,2199,2851,4349,5058,5079,7177,7959,8522,8886,10543,10832,10839,13359,13719,
99,215,2200,2852,4350,5059,5080,7178,7960,8523,8887,10544,10833,10840,13360,13720,
100,216,2201,2853,4351,5060,5081,7179,7961,8524,8888,10545,10834,10841,13361,13721,
101,217,2202,2854,4352,5061,5082,7180,7962,8525,8889,10546,10835,10842,13362,13722,
102,218,2203,2855,4353,5062,5083,7181,7963,8526,8890,10547,10836,10843,13363,13723,
103,219,2204,2856,4354,5063,5084,7182,7964,8527,8891,10548,10837,10844,13364,13724,
104,220,2205,2857,4355,5064,5085,7183,7965,8528,8892,10549,10838,10845,13365,13725,
105,221,2206,2858,4356,5065,5086,7184,7966,8529,8893,10550,10839,10846,13366,13726,
106,222,2207,2859,4357,5066,5087,7185,7967,8530,8894,10551,10840,10847,13367,13727,
107,223,2208,2860,4358,5067,5088,7186,7968,8531,8895,10552,10841,10848,13368,13728,
108,224,2209,2861,4359,5068,5089,7187,7969,8532,8896,10553,10842,10849,13369,13729,
109,225,2210,2862,4360,5069,5090,7188,7970,8533,8897,10554,10843,10850,13370,13730,
110,226,2211,2863,4361,5070,5091,7189,7971,8534,8898,10555,10844,10851,13371,13731,
111,227,2212,2864,4362,5071,5092,7190,7972,8535,8899,10556,10845,10852,13372,13732,
112,228,2213,2865,4363,5072,5093,7191,7973,8536,8900,10557,10846,10853,13373,13733,
113,229,2214,2866,4364,5073,5094,7192,7974,8537,8901,10558,10847,10854,13374,13734,
114,230,2215,2867,4365,5074,5095,7193,7975,8538,8902,10559,10848,10855,13375,13735,
115,231,2216,2868,4366,5075,5096,7194,7976,8539,8903,10560,10849,10856,13376,13736,
116,232,2217,2869,4367,5076,5097,7195,7977,8540,8904,10561,10850,10857,13377,13737,
117,233,2218,2870,4368,5077,5098,7196,7978,8541,8905,10562,10851,10858,13378,13738,
118,234,2219,2871,4369,5078,5099,7197,7979,8542,8906,10563,10852,10859,13379,13739,
119,235,2220,2872,4370,5079,5100,7198,7980,8543,8907,10564,10853,10860,13380,13740,
120,236,2221,2873,4371,5080,5101,7199,7981,8544,8908,10565,10854,10861,13381,13741,
121,237,2222,2874,4372,5081,5102,6840,7982,8545,8909,10566,10855,10862,13382,13742,
122,238,2223,2875,4373,5082,5103,6841,7983,8546,8910,10567,10856,10863,13383,13743,
123,239,2224,2876,4374,5083,5104,6842,7984,8547,8911,10568,10857,10864,13384,13744,
124,240,2225,2877,4375,5084,5105,6843,7985,8548,8912,10569,10858,10865,13385,13745,
125,241,2226,2878,4376,5085,5106,6844,7986,8549,8913,10570,10859,10866,13386,13746,
126,242,2227,2879,4377,5086,5107,6845,7987,8550,8914,10571,10860,10867,13387,13747,
127,243,2228,2520,4378,5087,5108,6846,7988,8551,8915,10572,10861,10868,13388,13748,
128,244,2229,2521,4379,5088,5109,6847,7989,8552,8916,10573,10862,10869,13389,13749,
129,245,2230,2522,4380,5089,5110,6848,7990,8553,8917,10574,10863,10870,13390,13750,
130,246,2231,2523,4381,5090,5111,6849,7991,8554,8918,10575,10864,10871,13391,13751,
131,247,2232,2524,4382,5091,5112,6850,7992,8555,8919,10576,10865,10872,13392,13752,
132,248,2233,2525,4383,5092,5113,6851,7993,8556,8920,10577,10866,10873,13393,13753,
133,249,2234,2526,4384,5093,5114,6852,7994,8557,8921,10578,10867,10874,13394,13754,
134,250,2235,2527,4385,5094,5115,6853,7995,8558,8922,10579,10868,10875,13395,13755,
135,251,2236,2528,4386,5095,5116,6854,7996,8559,8923,10580,10869,10876,13396,13756,
136,252,2237,2529,4387,5096,5117,6855,7997,8560,8924,10581,10870,10877,13397,13757,
137,253,2238,2530,4388,5097,5118,6856,7998,8561,8925,10582,10871,10878,13398,13758,
138,254,2239,2531,4389,5098,5119,6857,7999,8562,8926,10583,10872,10879,13399,13759,
139,255,2240,2532,4390,5099,5120,6858,8000,8563,8927,10584,10873,10880,13400,13760,
140,256,2241,2533,4391,5100,5121,6859,8001,8564,8928,10585,10874,10881,13401,13761,
141,257,2242,2534,4392,5101,5122,6860,8002,8565,8929,10586,10875,10882,13402,13762,
142,258,2243,2535,4393,5102,5123,6861,8003,8566,8930,10587,10876,10883,13403,13763,
143,259,2244,2536,4394,5103,5124,6862,8004,8567,8931,10588,10877,10884,13404,13764,
144,260,2245,2537,4395,5104,5125,6863,8005,8568,8932,10589,10878,10885,13405,13765,
145,261,2246,2538,4396,5105,5126,6864,8006,8569,8933,10590,10879,10886,13406,13766,
146,262,2247,2539,4397,5106,5127,6865,8007,8570,8934,10591,10880,10887,13407,13767,
147,263,2248,2540,4398,5107,5128,6866,8008,8571,8935,10592,10881,10888,13408,13768,
148,264,2249,2541,4399,5108,5129,6867,8009,8572,8936,10593,10882,10889,13409,13769,
149,265,2250,2542,4400,5109,5130,6868,8010,8573,8937,10594,10883,10890,13410,13770,
150,266,2251,2543,4401,5110,5131,6869,8011,8574,8938,10595,10884,10891,13411,13771,
151,267,2252,2544,4402,5111,5132,6870,8012,8575,8939,10596,10885,10892,13412,13772,
152,268,2253,2545,4403,5112,5133,6871,8013,8576,8940,10597,10886,10893,13413,13773,
153,269,2254,2546,4404,5113,5134,6872,8014,8577,8941,10598,10887,10894,13414,13774,
154,270,2255,2547,4405,5114,5135,6873,8015,8578,8942,10599,10888,10895,13415,13775,
155,271,2256,2548,4406,5115,5136,6874,8016,8579,8943,10600,10889,10896,13416,13776,
156,272,2257,2549,4407,5116,5137,6875,8017,8580,8944,10601,10890,10897,13417,13777,
157,273,2258,2550,4408,5117,5138,6876,8018,8581,8945,10602,10891,10898,13418,13778,
158,274,2259,2551,4409,5118,5139,6877,8019,8582,8946,10603,10892,10899,13419,13779,
159,275,2260,2552,4410,5119,5140,6878,8020,8583,8947,10604,10893,10900,13420,13780,
160,276,2261,2553,4411,5120,5141,6879,8021,8584,8948,10605,10894,10901,13421,13781,
161,277,2262,2554,4412,5121,5142,6880,8022,8585,8949,10606,10895,10902,13422,13782,
162,278,2263,2555,4413,5122,5143,6881,8023,8586,8950,10607,10896,10903,13423,13783,
163,279,2264,2556,4414,5123,5144,6882,8024,8587,8951,10608,10897,10904,13424,13784,
164,280,2265,2557,4415,5124,5145,6883,8025,8588,8952,10609,10898,10905,13425,13785,
165,281,2266,2558,4416,5125,5146,6884,8026,8589,8953,10610,10899,10906,13426,13786,
166,282,2267,2559,4417,5126,5147,6885,8027,8590,8954,10611,10900,10907,13427,13787,
167,283,2268,2560,4418,5127,5148,6886,8028,8591,8955,10612,10901,10908,13428,13788,
168,284,2269,2561,4419,5128,5149,6887,8029,8592,8956,10613,10902,10909,13429,13789,
169,285,2270,2562,4420,5129,5150,6888,8030,8593,8957,10614,10903,10910,13430,13790,
170,286,2271,2563,4421,5130,5151,6889,8031,8594,8958,10615,10904,10911,13431,13791,
171,287,2272,2564,4422,5131,5152,6890,8032,8595,8959,10616,10905,10912,13432,13792,
172,288,2273,2565,4423,5132,5153,6891,8033,8596,8960,10617,10906,10913,13433,13793,
173,289,2274,2566,4424,5133,5154,6892,8034,8597,8961,10618,10907,10914,13434,13794,
174,290,2275,2567,4425,5134,5155,6893,8035,8598,8962,10619,10908,10915,13435,13795,
175,291,2276,2568,4426,5135,5156,6894,8036,8599,8963,10620,10909,10916,13436,13796,
176,292,2277,2569,4427,5136,5157,6895,8037,8600,8964,10621,10910,10917,13437,13797,
177,293,2278,2570,4428,5137,5158,6896,8038,8601,8965,10622,10911,10918,13438,13798,
178,294,2279,2571,4429,5138,5159,6897,8039,8602,8966,10623,10912,10919,13439,13799,
179,295,2280,2572,4430,5139,5160,6898,8040,8603,8967,10624,10913,10920,13440,13800,
180,296,2281,2573,4431,5140,5161,6899,8041,8604,8968,10625,10914,10921,13441,13801,
181,297,2282,2574,4432,5141,5162,6900,8042,8605,8969,10626,10915,10922,13442,13802,
182,298,2283,2575,4433,5142,5163,6901,8043,8606,8970,10627,10916,10923,13443,13803,
183,299,2284,2576,4434,5143,5164,6902,8044,8607,8971,10628,10917,10924,13444,13804,
184,300,2285,2577,4435,5144,5165,6903,8045,8608,8972,10629,10918,10925,13445,13805,
185,301,2286,2578,4436,5145,5166,6904,8046,8609,8973,10630,10919,10926,13446,13806,
186,302,2287,2579,4437,5146,5167,6905,8047,8610,8974,10631,10920,10927,13447,13807,
187,303,2288,2580,4438,5147,5168,6906,8048,8611,8975,10632,10921,10928,13448,13808,
188,304,2289,2581,4439,5148,5169,6907,8049,8612,8976,10633,10922,10929,13449,13809,
189,305,2290,2582,4440,5149,5170,6908,8050,8613,8977,10634,10923,10930,13450,13810,
190,306,2291,2583,4441,5150,5171,6909,8051,8614,8978,10635,10924,10931,13451,13811,
191,307,2292,2584,4442,5151,5172,6910,8052,8615,8979,10636,10925,10932,13452,13812,
192,308,2293,2585,4443,5152,5173,6911,8053,8616,8980,10637,10926,10933,13453,13813,
193,309,2294,2586,4444,5153,5174,6912,8054,8617,8981,10638,10927,10934,13454,13814,
194,310,2295,2587,4445,5154,5175,6913,8055,8618,8982,10639,10928,10935,13455,13815,
195,311,2296,2588,4446,5155,5176,6914,8056,8619,8983,10640,10929,10936,13456,13816,
196,312,2297,2589,4447,5156,5177,6915,8057,8620,8984,10641,10930,10937,13457,13817,
197,313,2298,2590,4448,5157,5178,6916,8058,8621,8985,10642,10931,10938,13458,13818,
198,314,2299,2591,4449,5158,5179,6917,8059,8622,8986,10643,10932,10939,13459,13819,
199,315,2300,2592,4450,5159,5180,6918,8060,8623,8987,10644,10933,10940,13460,13820,
200,316,2301,2593,4451,5160,5181,6919,8061,8624,8988,10645,10934,10941,13461,13821,
201,317,2302,2594,4452,5161,5182,6920,8062,8625,8989,10646,10935,10942,13462,13822,
202,318,2303,2595,4453,5162,5183,6921,8063,8626,8990,10647,10936,10943,13463,13823,
203,319,2304,2596,4454,5163,5184,6922,8064,8627,8991,10648,10937,10944,13464,13824,
204,320,2305,2597,4455,5164,5185,6923,8065,8628,8992,10649,10938,10945,13465,13825,
205,321,2306,2598,4456,5165,5186,6924,8066,8629,8993,10650,10939,10946,13466,13826,
206,322,2307,2599,4457,5166,5187,6925,8067,8630,8994,10651,10940,10947,13467,13827,
207,323,2308,2600,4458,5167,5188,6926,8068,8631,8995,10652,10941,10948,13468,13828,
208,324,2309,2601,4459,5168,5189,6927,8069,8632,8996,10653,10942,10949,13469,13829,
209,325,2310,2602,4460,5169,5190,6928,8070,8633,8997,10654,10943,10950,13470,13830,
210,326,2311,2603,4461,5170,5191,6929,8071,8634,8998,10655,10944,10951,13471,13831,
211,327,2312,2604,4462,5171,5192,6930,8072,8635,8999,10656,10945,10952,13472,13832,
212,328,2313,2605,4463,5172,5193,6931,8073,8636,8640,10657,10946,10953,13473,13833,
213,329,2314,2606,4464,5173,5194,6932,8074,8637,8641,10658,10947,10954,13474,13834,
214,330,2315,2607,4465,5174,5195,6933,8075,8638,8642,10659,10948,10955,13475,13835,
215,331,2316,2608,4466,5175,5196,6934,8076,8639,8643,10660,10949,10956,13476,13836,
216,332,2317,2609,4467,5176,5197,6935,8077,8280,8644,10661,10950,10957,13477,13837,
217,333,2318,2610,4468,5177,5198,6936,8078,8281,8645,10662,10951,10958,13478,13838,
218,334,2319,2611,4469,5178,5199,6937,8079,8282,8646,10663,10952,10959,13479,13839,
219,335,2320,2612,4470,5179,5200,6938,8080,8283,8647,10664,10953,10960,13480,13840,
220,336,2321,2613,4471,5180,5201,6939,8081,8284,8648,10665,10954,10961,13481,13841,
221,337,2322,2614,4472,5181,5202,6940,8082,8285,8649,10666,10955,10962,13482,13842,
222,338,2323,2615,4473,5182,5203,6941,8083,8286,8650,10667,10956,10963,13483,13843,
223,339,2324,2616,4474,5183,5204,6942,8084,8287,8651,10668,10957,10964,13484,13844,
224,340,2325,2617,4475,5184,5205,6943,8085,8288,8652,10669,10958,10965,13485,13845,
225,341,2326,2618,4476,5185,5206,6944,8086,8289,8653,10670,10959,10966,13486,13846,
226,342,2327,2619,4477,5186,5207,6945,8087,8290,8654,10671,10960,10967,13487,13847,
227,343,2328,2620,4478,5187,5208,6946,8088,8291,8655,10672,10961,10968,13488,13848,
228,344,2329,2621,4479,5188,5209,6947,8089,8292,8656,10673,10962,10969,13489,13849,
229,345,2330,2622,4480,5189,5210,6948,8090,8293,8657,10674,10963,10970,13490,13850,
230,346,2331,2623,4481,5190,5211,6949,8091,8294,8658,10675,10964,10971,13491,13851,
231,347,2332,2624,4482,5191,5212,6950,8092,8295,8659,10676,10965,10972,13492,13852,
232,348,2333,2625,4483,5192,5213,6951,8093,8296,8660,10677,10966,10973,13493,13853,
233,349,2334,2626,4484,5193,5214,6952,8094,8297,8661,10678,10967,10974,13494,13854,
234,350,2335,2627,4485,5194,5215,6953,8095,8298,8662,10679,10968,10975,13495,13855,
235,351,2336,2628,4486,5195,5216,6954,8096,8299,8663,10680,10969,10976,13496,13856,
236,352,2337,2629,4487,5196,5217,6955,8097,8300,8664,10681,10970,10977,13497,13857,
237,353,2338,2630,4488,5197,5218,6956,8098,8301,8665,10682,10971,10978,13498,13858,
238,354,2339,2631,4489,5198,5219,6957,8099,8302,8666,10683,10972,10979,13499,13859,
239,355,2340,2632,4490,5199,5220,6958,8100,8303,8667,10684,10973,10980,13500,13860,
240,356,2341,2633,4491,5200,5221,6959,8101,8304,8668,10685,10974,10981,13501,13861,
241,357,2342,2634,4492,5201,5222,6960,8102,8305,8669,10686,10975,10982,13502,13862,
242,358,2343,2635,4493,5202,5223,6961,8103,8306,8670,10687,10976,10983,13503,13863,
243,359,2344,2636,4494,5203,5224,6962,8104,8307,8671,10688,10977,10984,13504,13864,
0,244,2345,2637,4495,5204,5225,6963,8105,8308,8672,10689,10978,10985,13505,13865,
1,245,2346,2638,4496,5205,5226,6964,8106,8309,8673,10690,10979,10986,13506,13866,
2,246,2347,2639,4497,5206,5227,6965,8107,8310,8674,10691,10980,10987,13507,13867,
3,247,2348,2640,4498,5207,5228,6966,8108,8311,8675,10692,10981,10988,13508,13868,
4,248,2349,2641,4499,5208,5229,6967,8109,8312,8676,10693,10982,10989,13509,13869,
5,249,2350,2642,4500,5209,5230,6968,8110,8313,8677,10694,10983,10990,13510,13870,
6,250,2351,2643,4501,5210,5231,6969,8111,8314,8678,10695,10984,10991,13511,13871,
7,251,2352,2644,4502,5211,5232,6970,8112,8315,8679,10696,10985,10992,13512,13872,
8,252,2353,2645,4503,5212,5233,6971,8113,8316,8680,10697,10986,10993,13513,13873,
9,253,2354,2646,4504,5213,5234,6972,8114,8317,8681,10698,10987,10994,13514,13874,
10,254,2355,2647,4505,5214,5235,6973,8115,8318,8682,10699,10988,10995,13515,13875,
11,255,2356,2648,4506,5215,5236,6974,8116,8319,8683,10700,10989,10996,13516,13876,
12,256,2357,2649,4507,5216,5237,6975,8117,8320,8684,10701,10990,10997,13517,13877,
13,257,2358,2650,4508,5217,5238,6976,8118,8321,8685,10702,10991,10998,13518,13878,
14,258,2359,2651,4509,5218,5239,6977,8119,8322,8686,10703,10992,10999,13519,13879,
15,259,2360,2652,4510,5219,5240,6978,8120,8323,8687,10704,10993,11000,13520,13880,
16,260,2361,2653,4511,5220,5241,6979,8121,8324,8688,10705,10994,11001,13521,13881,
17,261,2362,2654,4512,5221,5242,6980,8122,8325,8689,10706,10995,11002,13522,13882,
18,262,2363,2655,4513,5222,5243,6981,8123,8326,8690,10707,10996,11003,13523,13883,
19,263,2364,2656,4514,5223,5244,6982,8124,8327,8691,10708,10997,11004,13524,13884,
20,264,2365,2657,4515,5224,5245,6983,8125,8328,8692,10709,10998,11005,13525,13885,
21,265,2366,2658,4516,5225,5246,6984,8126,8329,8693,10710,10999,11006,13526,13886,
22,266,2367,2659,4517,5226,5247,6985,8127,8330,8694,10711,11000,11007,13527,13887,
23,267,2368,2660,4518,5227,5248,6986,8128,8331,8695,10712,11001,11008,13528,13888,
24,268,2369,2661,4519,5228,5249,6987,8129,8332,8696,10713,11002,11009,13529,13889,
25,269,2370,2662,4520,5229,5250,6988,8130,8333,8697,10714,11003,11010,13530,13890,
26,270,2371,2663,4521,5230,5251,6989,8131,8334,8698,10715,11004,11011,13531,13891,
27,271,2372,2664,4522,5231,5252,6990,8132,8335,8699,10716,11005,11012,13532,13892,
28,272,2373,2665,4523,5232,5253,6991,8133,8336,8700,10717,11006,11013,13533,13893,
29,273,2374,2666,4524,5233,5254,6992,8134,8337,8701,10718,11007,11014,13534,13894,
30,274,2375,2667,4525,5234,5255,6993,8135,8338,8702,10719,11008,11015,13535,13895,
31,275,2376,2668,4526,5235,5256,6994,8136,8339,8703,10720,11009,11016,13536,13896,
32,276,2377,2669,4527,5236,5257,6995,8137,8340,8704,10721,11010,11017,13537,13897,
33,277,2378,2670,4528,5237,5258,6996,8138,8341,8705,10722,11011,11018,13538,13898,
34,278,2379,2671,4529,5238,5259,6997,8139,8342,8706,10723,11012,11019,13539,13899,
35,279,2380,2672,4530,5239,5260,6998,8140,8343,8707,10724,11013,11020,13540,13900,
36,280,2381,2673,4531,5240,5261,6999,8141,8344,8708,10725,11014,11021,13541,13901,
37,281,2382,2674,4532,5241,5262,7000,8142,8345,8709,10726,11015,11022,13542,13902,
38,282,2383,2675,4533,5242,5263,7001,8143,8346,8710,10727,11016,11023,13543,13903,
39,283,2384,2676,4534,5243,5264,7002,8144,8347,8711,10728,11017,11024,13544,13904,
40,284,2385,2677,4535,5244,5265,7003,8145,8348,8712,10729,11018,11025,13545,13905,
41,285,2386,2678,4536,5245,5266,7004,8146,8349,8713,10730,11019,11026,13546,13906,
42,286,2387,2679,4537,5246,5267,7005,8147,8350,8714,10731,11020,11027,13547,13907,
43,287,2388,2680,4538,5247,5268,7006,8148,8351,8715,10732,11021,11028,13548,13908,
44,288,2389,2681,4539,5248,5269,7007,8149,8352,8716,10733,11022,11029,13549,13909,
45,289,2390,2682,4540,5249,5270,7008,8150,8353,8717,10734,11023,11030,13550,13910,
46,290,2391,2683,4541,5250,5271,7009,8151,8354,8718,10735,11024,11031,13551,13911,
47,291,2392,2684,4542,5251,5272,7010,8152,8355,8719,10736,11025,11032,13552,13912,
48,292,2393,2685,4543,5252,5273,7011,8153,8356,8720,10737,11026,11033,13553,13913,
49,293,2394,2686,4544,5253,5274,7012,8154,8357,8721,10738,11027,11034,13554,13914,
50,294,2395,2687,4545,5254,5275,7013,8155,8358,8722,10739,11028,11035,13555,13915,
51,295,2396,2688,4546,5255,5276,7014,8156,8359,8723,10740,11029,11036,13556,13916,
52,296,2397,2689,4547,5256,5277,7015,8157,8360,8724,10741,11030,11037,13557,13917,
53,297,2398,2690,4548,5257,5278,7016,8158,8361,8725,10742,11031,11038,13558,13918,
54,298,2399,2691,4549,5258,5279,7017,8159,8362,8726,10743,11032,11039,13559,13919,
55,299,2400,2692,4550,5259,5280,7018,8160,8363,8727,10744,11033,11040,13560,13920,
56,300,2401,2693,4551,5260,5281,7019,8161,8364,8728,10745,11034,11041,13561,13921,
57,301,2402,2694,4552,5261,5282,7020,8162,8365,8729,10746,11035,11042,13562,13922,
58,302,2403,2695,4553,5262,5283,7021,8163,8366,8730,10747,11036,11043,13563,13923,
59,303,2404,2696,4554,5263,5284,7022,8164,8367,8731,10748,11037,11044,13564,13924,
60,304,2405,2697,4555,5264,5285,7023,8165,8368,8732,10749,11038,11045,13565,13925,
61,305,2406,2698,4556,5265,5286,7024,8166,8369,8733,10750,11039,11046,13566,13926,
62,306,2407,2699,4557,5266,5287,7025,8167,8370,8734,10751,11040,11047,13567,13927,
63,307,2408,2700,4558,5267,5288,7026,8168,8371,8735,10752,11041,11048,13568,13928,
64,308,2409,2701,4559,5268,5289,7027,8169,8372,8736,10753,11042,11049,13569,13929,
65,309,2410,2702,4560,5269,5290,7028,8170,8373,8737,10754,11043,11050,13570,13930,
66,310,2411,2703,4561,5270,5291,7029,8171,8374,8738,10755,11044,11051,13571,13931,
67,311,2412,2704,4562,5271,5292,7030,8172,8375,8739,10756,11045,11052,13572,13932,
68,312,2413,2705,4563,5272,5293,7031,8173,8376,8740,10757,11046,11053,13573,13933,
69,313,2414,2706,4564,5273,5294,7032,8174,8377,8741,10758,11047,11054,13574,13934,
70,314,2415,2707,4565,5274,5295,7033,8175,8378,8742,10759,11048,11055,13575,13935,
71,315,2416,2708,4566,5275,5296,7034,8176,8379,8743,10760,11049,11056,13576,13936,
72,316,2417,2709,4567,5276,5297,7035,8177,8380,8744,10761,11050,11057,13577,13937,
73,317,2418,2710,4568,5277,5298,7036,8178,8381,8745,10762,11051,11058,13578,13938,
74,318,2419,2711,4569,5278,5299,7037,8179,8382,8746,10763,11052,11059,13579,13939,
75,319,2420,2712,4570,5279,5300,7038,8180,8383,8747,10764,11053,11060,13580,13940,
76,320,2421,2713,4571,5280,5301,7039,8181,8384,8748,10765,11054,11061,13581,13941,
77,321,2422,2714,4572,5281,5302,7040,8182,8385,8749,10766,11055,11062,13582,13942,
78,322,2423,2715,4573,5282,5303,7041,8183,8386,8750,10767,11056,11063,13583,13943,
79,323,2424,2716,4574,5283,5304,7042,8184,8387,8751,10768,11057,11064,13584,13944,
80,324,2425,2717,4575,5284,5305,7043,8185,8388,8752,10769,11058,11065,13585,13945,
81,325,2426,2718,4576,5285,5306,7044,8186,8389,8753,10770,11059,11066,13586,13946,
82,326,2427,2719,4577,5286,5307,7045,8187,8390,8754,10771,11060,11067,13587,13947,
83,327,2428,2720,4578,5287,5308,7046,8188,8391,8755,10772,11061,11068,13588,13948,
84,328,2429,2721,4579,5288,5309,7047,8189,8392,8756,10773,11062,11069,13589,13949,
85,329,2430,2722,4580,5289,5310,7048,8190,8393,8757,10774,11063,11070,13590,13950,
86,330,2431,2723,4581,5290,5311,7049,8191,8394,8758,10775,11064,11071,13591,13951,
87,331,2432,2724,4582,5291,5312,7050,8192,8395,8759,10776,11065,11072,13592,13952,
88,332,2433,2725,4583,5292,5313,7051,8193,8396,8760,10777,11066,11073,13593,13953,
89,333,2434,2726,4584,5293,5314,7052,8194,8397,8761,10778,11067,11074,13594,13954,
90,334,2435,2727,4585,5294,5315,7053,8195,8398,8762,10779,11068,11075,13595,13955,
91,335,2436,2728,4586,5295,5316,7054,8196,8399,8763,10780,11069,11076,13596,13956,
92,336,2437,2729,4587,5296,5317,7055,8197,8400,8764,10781,11070,11077,13597,13957,
93,337,2438,2730,4588,5297,5318,7056,8198,8401,8765,10782,11071,11078,13598,13958,
94,338,2439,2731,4589,5298,5319,7057,8199,8402,8766,10783,11072,11079,13599,13959,
95,339,2440,2732,4590,5299,5320,7058,8200,8403,8767,10784,11073,11080,13600,13960,
96,340,2441,2733,4591,5300,5321,7059,8201,8404,8768,10785,11074,11081,13601,13961,
97,341,2442,2734,4592,5301,5322,7060,8202,8405,8769,10786,11075,11082,13602,13962,
98,342,2443,2735,4593,5302,5323,7061,8203,8406,8770,10787,11076,11083,13603,13963,
99,343,2444,2736,4594,5303,5324,7062,8204,8407,8771,10788,11077,11084,13604,13964,
100,344,2445,2737,4595,5304,5325,7063,8205,8408,8772,10789,11078,11085,13605,13965,
101,345,2446,2738,4596,5305,5326,7064,8206,8409,8773,10790,11079,11086,13606,13966,
102,346,2447,2739,4597,5306,5327,7065,8207,8410,8774,10791,11080,11087,13607,13967,
103,347,2448,2740,4598,5307,5328,7066,8208,8411,8775,10792,11081,11088,13608,13968,
104,348,2449,2741,4599,5308,5329,7067,8209,8412,8776,10793,11082,11089,13609,13969,
105,349,2450,2742,4600,5309,5330,7068,8210,8413,8777,10794,11083,11090,13610,13970,
106,350,2451,2743,4601,5310,5331,7069,8211,8414,8778,10795,11084,11091,13611,13971,
107,351,2452,2744,4602,5311,5332,7070,8212,8415,8779,10796,11085,11092,13612,13972,
108,352,2453,2745,4603,5312,5333,7071,8213,8416,8780,10797,11086,11093,13613,13973,
109,353,2454,2746,4604,5313,5334,7072,8214,8417,8781,10798,11087,11094,13614,13974,
110,354,2455,2747,4605,5314,5335,7073,8215,8418,8782,10799,11088,11095,13615,13975,
111,355,2456,2748,4606,5315,5336,7074,8216,8419,8783,10440,11089,11096,13616,13976,
112,356,2457,2749,4607,5316,5337,7075,8217,8420,8784,10441,11090,11097,13617,13977,
113,357,2458,2750,4608,5317,5338,7076,8218,8421,8785,10442,11091,11098,13618,13978,
114,358,2459,2751,4609,5318,5339,7077,8219,8422,8786,10443,11092,11099,13619,13979,
115,359,2460,2752,4610,5319,5340,7078,8220,8423,8787,10444,11093,11100,13620,13980,
0,116,2461,2753,4611,5320,5341,7079,8221,8424,8788,10445,11094,11101,13621,13981,
1,117,2462,2754,4612,5321,5342,7080,8222,8425,8789,10446,11095,11102,13622,13982,
2,118,2463,2755,4613,5322,5343,7081,8223,8426,8790,10447,11096,11103,13623,13983,
3,119,2464,2756,4614,5323,5344,7082,8224,8427,8791,10448,11097,11104,13624,13984,
4,120,2465,2757,4615,5324,5345,7083,8225,8428,8792,10449,11098,11105,13625,13985,
5,121,2466,2758,4616,5325,5346,7084,8226,8429,8793,10450,11099,11106,13626,13986,
6,122,2467,2759,4617,5326,5347,7085,8227,8430,8794,10451,11100,11107,13627,13987,
7,123,2468,2760,4618,5327,5348,7086,8228,8431,8795,10452,11101,11108,13628,13988,
8,124,2469,2761,4619,5328,5349,7087,8229,8432,8796,10453,11102,11109,13629,13989,
9,125,2470,2762,4620,5329,5350,7088,8230,8433,8797,10454,11103,11110,13630,13990,
10,126,2471,2763,4621,5330,5351,7089,8231,8434,8798,10455,11104,11111,13631,13991,
11,127,2472,2764,4622,5331,5352,7090,8232,8435,8799,10456,11105,11112,13632,13992,
12,128,2473,2765,4623,5332,5353,7091,8233,8436,8800,10457,11106,11113,13633,13993,
13,129,2474,2766,4624,5333,5354,7092,8234,8437,8801,10458,11107,11114,13634,13994,
14,130,2475,2767,4625,5334,5355,7093,8235,8438,8802,10459,11108,11115,13635,13995,
15,131,2476,2768,4626,5335,5356,7094,8236,8439,8803,10460,11109,11116,13636,13996,
16,132,2477,2769,4627,5336,5357,7095,8237,8440,8804,10461,11110,11117,13637,13997,
17,133,2478,2770,4628,5337,5358,7096,8238,8441,8805,10462,11111,11118,13638,13998,
18,134,2479,2771,4629,5338,5359,7097,8239,8442,8806,10463,11112,11119,13639,13999,
19,135,2480,2772,4630,5339,5360,7098,8240,8443,8807,10464,11113,11120,13640,14000,
20,136,2481,2773,4631,5340,5361,7099,8241,8444,8808,10465,11114,11121,13641,14001,
21,137,2482,2774,4632,5341,5362,7100,8242,8445,8809,10466,11115,11122,13642,14002,
22,138,2483,2775,4633,5342,5363,7101,8243,8446,8810,10467,11116,11123,13643,14003,
23,139,2484,2776,4634,5343,5364,7102,8244,8447,8811,10468,11117,11124,13644,14004,
24,140,2485,2777,4635,5344,5365,7103,8245,8448,8812,10469,11118,11125,13645,14005,
25,141,2486,2778,4636,5345,5366,7104,8246,8449,8813,10470,11119,11126,13646,14006,
26,142,2487,2779,4637,5346,5367,7105,8247,8450,8814,10471,11120,11127,13647,14007,
27,143,2488,2780,4638,5347,5368,7106,8248,8451,8815,10472,11121,11128,13648,14008,
28,144,2489,2781,4639,5348,5369,7107,8249,8452,8816,10473,11122,11129,13649,14009,
29,145,2490,2782,4640,5349,5370,7108,8250,8453,8817,10474,11123,11130,13650,14010,
30,146,2491,2783,4641,5350,5371,7109,8251,8454,8818,10475,11124,11131,13651,14011,
31,147,2492,2784,4642,5351,5372,7110,8252,8455,8819,10476,11125,11132,13652,14012,
32,148,2493,2785,4643,5352,5373,7111,8253,8456,8820,10477,11126,11133,13653,14013,
33,149,2494,2786,4644,5353,5374,7112,8254,8457,8821,10478,11127,11134,13654,14014,
34,150,2495,2787,4645,5354,5375,7113,8255,8458,8822,10479,11128,11135,13655,14015,
35,151,2496,2788,4646,5355,5376,7114,8256,8459,8823,10480,11129,11136,13656,14016,
36,152,2497,2789,4647,5356,5377,7115,8257,8460,8824,10481,11130,11137,13657,14017,
37,153,2498,2790,4648,5357,5378,7116,8258,8461,8825,10482,11131,11138,13658,14018,
38,154,2499,2791,4649,5358,5379,7117,8259,8462,8826,10483,11132,11139,13659,14019,
39,155,2500,2792,4650,5359,5380,7118,8260,8463,8827,10484,11133,11140,13660,14020,
40,156,2501,2793,4651,5360,5381,7119,8261,8464,8828,10485,11134,11141,13661,14021,
41,157,2502,2794,4652,5361,5382,7120,8262,8465,8829,10486,11135,11142,13662,14022,
42,158,2503,2795,4653,5362,5383,7121,8263,8466,8830,10487,11136,11143,13663,14023,
43,159,2504,2796,4654,5363,5384,7122,8264,8467,8831,10488,11137,11144,13664,14024,
44,160,2505,2797,4655,5364,5385,7123,8265,8468,8832,10489,11138,11145,13665,14025,
45,161,2506,2798,4656,5365,5386,7124,8266,8469,8833,10490,11139,11146,13666,14026,
46,162,2507,2799,4657,5366,5387,7125,8267,8470,8834,10491,11140,11147,13667,14027,
47,163,2508,2800,4658,5367,5388,7126,8268,8471,8835,10492,11141,11148,13668,14028,
48,164,2509,2801,4659,5368,5389,7127,8269,8472,8836,10493,11142,11149,13669,14029,
49,165,2510,2802,4660,5369,5390,7128,8270,8473,8837,10494,11143,11150,13670,14030,
50,166,2511,2803,4661,5370,5391,7129,8271,8474,8838,10495,11144,11151,13671,14031,
51,167,2512,2804,4662,5371,5392,7130,8272,8475,8839,10496,11145,11152,13672,14032,
52,168,2513,2805,4663,5372,5393,7131,8273,8476,8840,10497,11146,11153,13673,14033,
53,169,2514,2806,4664,5373,5394,7132,8274,8477,8841,10498,11147,11154,13674,14034,
54,170,2515,2807,4665,5374,5395,7133,8275,8478,8842,10499,11148,11155,13675,14035,
55,171,2516,2808,4666,5375,5396,7134,8276,8479,8843,10500,11149,11156,13676,14036,
56,172,2517,2809,4667,5376,5397,7135,8277,8480,8844,10501,11150,11157,13677,14037,
57,173,2518,2810,4668,5377,5398,7136,8278,8481,8845,10502,11151,11158,13678,14038,
58,174,2519,2811,4669,5378,5399,7137,8279,8482,8846,10503,11152,11159,13679,14039,
1176,1335,2520,3318,4306,5400,5881,6299,7610,8280,8433,11160,11389,12023,13680,14040,
1177,1336,2521,3319,4307,5401,5882,6300,7611,8281,8434,11161,11390,12024,13681,14041,
1178,1337,2522,3320,4308,5402,5883,6301,7612,8282,8435,11162,11391,12025,13682,14042,
1179,1338,2523,3321,4309,5403,5884,6302,7613,8283,8436,11163,11392,12026,13683,14043,
1180,1339,2524,3322,4310,5404,5885,6303,7614,8284,8437,11164,11393,12027,13684,14044,
1181,1340,2525,3323,4311,5405,5886,6304,7615,8285,8438,11165,11394,12028,13685,14045,
1182,1341,2526,3324,4312,5406,5887,6305,7616,8286,8439,11166,11395,12029,13686,14046,
1183,1342,2527,3325,4313,5407,5888,6306,7617,8287,8440,11167,11396,12030,13687,14047,
1184,1343,2528,3326,4314,5408,5889,6307,7618,8288,8441,11168,11397,12031,13688,14048,
1185,1344,2529,3327,4315,5409,5890,6308,7619,8289,8442,11169,11398,12032,13689,14049,
1186,1345,2530,3328,4316,5410,5891,6309,7620,8290,8443,11170,11399,12033,13690,14050,
1187,1346,2531,3329,4317,5411,5892,6310,7621,8291,8444,11171,11400,12034,13691,14051,
1188,1347,2532,3330,4318,5412,5893,6311,7622,8292,8445,11172,11401,12035,13692,14052,
1189,1348,2533,3331,4319,5413,5894,6312,7623,8293,8446,11173,11402,12036,13693,14053,
1190,1349,2534,3332,3960,5414,5895,6313,7624,8294,8447,11174,11403,12037,13694,14054,
1191,1350,2535,3333,3961,5415,5896,6314,7625,8295,8448,11175,11404,12038,13695,14055,
1192,1351,2536,3334,3962,5416,5897,6315,7626,8296,8449,11176,11405,12039,13696,14056,
1193,1352,2537,3335,3963,5417,5898,6316,7627,8297,8450,11177,11406,12040,13697,14057,
1194,1353,2538,3336,3964,5418,5899,6317,7628,8298,8451,11178,11407,12041,13698,14058,
1195,1354,2539,3337,3965,5419,5900,6318,7629,8299,8452,11179,11408,12042,13699,14059,
1196,1355,2540,3338,3966,5420,5901,6319,7630,8300,8453,11180,11409,12043,13700,14060,
1197,1356,2541,3339,3967,5421,5902,6320,7631,8301,8454,11181,11410,12044,13701,14061,
1198,1357,2542,3340,3968,5422,5903,6321,7632,8302,8455,11182,11411,12045,13702,14062,
1199,1358,2543,3341,3969,5423,5904,6322,7633,8303,8456,11183,11412,12046,13703,14063,
1200,1359,2544,3342,3970,5424,5905,6323,7634,8304,8457,11184,11413,12047,13704,14064,
1201,1360,2545,3343,3971,5425,5906,6324,7635,8305,8458,11185,11414,12048,13705,14065,
1202,1361,2546,3344,3972,5426,5907,6325,7636,8306,8459,11186,11415,12049,13706,14066,
1203,1362,2547,3345,3973,5427,5908,6326,7637,8307,8460,11187,11416,12050,13707,14067,
1204,1363,2548,3346,3974,5428,5909,6327,7638,8308,8461,11188,11417,12051,13708,14068,
1205,1364,2549,3347,3975,5429,5910,6328,7639,8309,8462,11189,11418,12052,13709,14069,
1206,1365,2550,3348,3976,5430,5911,6329,7640,8310,8463,11190,11419,12053,13710,14070,
1207,1366,2551,3349,3977,5431,5912,6330,7641,8311,8464,11191,11420,12054,13711,14071,
1208,1367,2552,3350,3978,5432,5913,6331,7642,8312,8465,11192,11421,12055,13712,14072,
1209,1368,2553,3351,3979,5433,5914,6332,7643,8313,8466,11193,11422,12056,13713,14073,
1210,1369,2554,3352,3980,5434,5915,6333,7644,8314,8467,11194,11423,12057,13714,14074,
1211,1370,2555,3353,3981,5435,5916,6334,7645,8315,8468,11195,11424,12058,13715,14075,
1212,1371,2556,3354,3982,5436,5917,6335,7646,8316,8469,11196,11425,12059,13716,14076,
1213,1372,2557,3355,3983,5437,5918,6336,7647,8317,8470,11197,11426,12060,13717,14077,
1214,1373,2558,3356,3984,5438,5919,6337,7648,8318,8471,11198,11427,12061,13718,14078,
1215,1374,2559,3357,3985,5439,5920,6338,7649,8319,8472,11199,11428,12062,13719,14079,
1216,1375,2560,3358,3986,5440,5921,6339,7650,8320,8473,11200,11429,12063,13720,14080,
1217,1376,2561,3359,3987,5441,5922,6340,7651,8321,8474,11201,11430,12064,13721,14081,
1218,1377,2562,3360,3988,5442,5923,6341,7652,8322,8475,11202,11431,12065,13722,14082,
1219,1378,2563,3361,3989,5443,5924,6342,7653,8323,8476,11203,11432,12066,13723,14083,
1220,1379,2564,3362,3990,5444,5925,6343,7654,8324,8477,11204,11433,12067,13724,14084,
1221,1380,2565,3363,3991,5445,5926,6344,7655,8325,8478,11205,11434,12068,13725,14085,
1222,1381,2566,3364,3992,5446,5927,6345,7656,8326,8479,11206,11435,12069,13726,14086,
1223,1382,2567,3365,3993,5447,5928,6346,7657,8327,8480,11207,11436,12070,13727,14087,
1224,1383,2568,3366,3994,5448,5929,6347,7658,8328,8481,11208,11437,12071,13728,14088,
1225,1384,2569,3367,3995,5449,5930,6348,7659,8329,8482,11209,11438,12072,13729,14089,
1226,1385,2570,3368,3996,5450,5931,6349,7660,8330,8483,11210,11439,12073,13730,14090,
1227,1386,2571,3369,3997,5451,5932,6350,7661,8331,8484,11211,11440,12074,13731,14091,
1228,1387,2572,3370,3998,5452,5933,6351,7662,8332,8485,11212,11441,12075,13732,14092,
1229,1388,2573,3371,3999,5453,5934,6352,7663,8333,8486,11213,11442,12076,13733,14093,
1230,1389,2574,3372,4000,5454,5935,6353,7664,8334,8487,11214,11443,12077,13734,14094,
1231,1390,2575,3373,4001,5455,5936,6354,7665,8335,8488,11215,11444,12078,13735,14095,
1232,1391,2576,3374,4002,5456,5937,6355,7666,8336,8489,11216,11445,12079,13736,14096,
1233,1392,2577,3375,4003,5457,5938,6356,7667,8337,8490,11217,11446,12080,13737,14097,
1234,1393,2578,3376,4004,5458,5939,6357,7668,8338,8491,11218,11447,12081,13738,14098,
1235,1394,2579,3377,4005,5459,5940,6358,7669,8339,8492,11219,11448,12082,13739,14099,
1236,1395,2580,3378,4006,5460,5941,6359,7670,8340,8493,11220,11449,12083,13740,14100,
1237,1396,2581,3379,4007,5461,5942,6360,7671,8341,8494,11221,11450,12084,13741,14101,
1238,1397,2582,3380,4008,5462,5943,6361,7672,8342,8495,11222,11451,12085,13742,14102,
1239,1398,2583,3381,4009,5463,5944,6362,7673,8343,8496,11223,11452,12086,13743,14103,
1240,1399,2584,3382,4010,5464,5945,6363,7674,8344,8497,11224,11453,12087,13744,14104,
1241,1400,2585,3383,4011,5465,5946,6364,7675,8345,8498,11225,11454,12088,13745,14105,
1242,1401,2586,3384,4012,5466,5947,6365,7676,8346,8499,11226,11455,12089,13746,14106,
1243,1402,2587,3385,4013,5467,5948,6366,7677,8347,8500,11227,11456,12090,13747,14107,
1244,1403,2588,3386,4014,5468,5949,6367,7678,8348,8501,11228,11457,12091,13748,14108,
1245,1404,2589,3387,4015,5469,5950,6368,7679,8349,8502,11229,11458,12092,13749,14109,
1246,1405,2590,3388,4016,5470,5951,6369,7680,8350,8503,11230,11459,12093,13750,14110,
1247,1406,2591,3389,4017,5471,5952,6370,7681,8351,8504,11231,11460,12094,13751,14111,
1248,1407,2592,3390,4018,5472,5953,6371,7682,8352,8505,11232,11461,12095,13752,14112,
1249,1408,2593,3391,4019,5473,5954,6372,7683,8353,8506,11233,11462,12096,13753,14113,
1250,1409,2594,3392,4020,5474,5955,6373,7684,8354,8507,11234,11463,12097,13754,14114,
1251,1410,2595,3393,4021,5475,5956,6374,7685,8355,8508,11235,11464,12098,13755,14115,
1252,1411,2596,3394,4022,5476,5957,6375,7686,8356,8509,11236,11465,12099,13756,14116,
1253,1412,2597,3395,4023,5477,5958,6376,7687,8357,8510,11237,11466,12100,13757,14117,
1254,1413,2598,3396,4024,5478,5959,6377,7688,8358,8511,11238,11467,12101,13758,14118,
1255,1414,2599,3397,4025,5479,5960,6378,7689,8359,8512,11239,11468,12102,13759,14119,
1256,1415,2600,3398,4026,5480,5961,6379,7690,8360,8513,11240,11469,12103,13760,14120,
1257,1416,2601,3399,4027,5481,5962,6380,7691,8361,8514,11241,11470,12104,13761,14121,
1258,1417,2602,3400,4028,5482,5963,6381,7692,8362,8515,11242,11471,12105,13762,14122,
1259,1418,2603,3401,4029,5483,5964,6382,7693,8363,8516,11243,11472,12106,13763,14123,
1260,1419,2604,3402,4030,5484,5965,6383,7694,8364,8517,11244,11473,12107,13764,14124,
1261,1420,2605,3403,4031,5485,5966,6384,7695,8365,8518,11245,11474,12108,13765,14125,
1262,1421,2606,3404,4032,5486,5967,6385,7696,8366,8519,11246,11475,12109,13766,14126,
1263,1422,2607,3405,4033,5487,5968,6386,7697,8367,8520,11247,11476,12110,13767,14127,
1264,1423,2608,3406,4034,5488,5969,6387,7698,8368,8521,11248,11477,12111,13768,14128,
1265,1424,2609,3407,4035,5489,5970,6388,7699,8369,8522,11249,11478,12112,13769,14129,
1266,1425,2610,3408,4036,5490,5971,6389,7700,8370,8523,11250,11479,12113,13770,14130,
1267,1426,2611,3409,4037,5491,5972,6390,7701,8371,8524,11251,11480,12114,13771,14131,
1268,1427,2612,3410,4038,5492,5973,6391,7702,8372,8525,11252,11481,12115,13772,14132,
1269,1428,2613,3411,4039,5493,5974,6392,7703,8373,8526,11253,11482,12116,13773,14133,
1270,1429,2614,3412,4040,5494,5975,6393,7704,8374,8527,11254,11483,12117,13774,14134,
1271,1430,2615,3413,4041,5495,5976,6394,7705,8375,8528,11255,11484,12118,13775,14135,
1272,1431,2616,3414,4042,5496,5977,6395,7706,8376,8529,11256,11485,12119,13776,14136,
1273,1432,2617,3415,4043,5497,5978,6396,7707,8377,8530,11257,11486,12120,13777,14137,
1274,1433,2618,3416,4044,5498,5979,6397,7708,8378,8531,11258,11487,12121,13778,14138,
1275,1434,2619,3417,4045,5499,5980,6398,7709,8379,8532,11259,11488,12122,13779,14139,
1276,1435,2620,3418,4046,5500,5981,6399,7710,8380,8533,11260,11489,12123,13780,14140,
1277,1436,2621,3419,4047,5501,5982,6400,7711,8381,8534,11261,11490,12124,13781,14141,
1278,1437,2622,3420,4048,5502,5983,6401,7712,8382,8535,11262,11491,12125,13782,14142,
1279,1438,2623,3421,4049,5503,5984,6402,7713,8383,8536,11263,11492,12126,13783,14143,
1280,1439,2624,3422,4050,5504,5985,6403,7714,8384,8537,11264,11493,12127,13784,14144,
1080,1281,2625,3423,4051,5505,5986,6404,7715,8385,8538,11265,11494,12128,13785,14145,
1081,1282,2626,3424,4052,5506,5987,6405,7716,8386,8539,11266,11495,12129,13786,14146,
1082,1283,2627,3425,4053,5507,5988,6406,7717,8387,8540,11267,11496,12130,13787,14147,
1083,1284,2628,3426,4054,5508,5989,6407,7718,8388,8541,11268,11497,12131,13788,14148,
1084,1285,2629,3427,4055,5509,5990,6408,7719,8389,8542,11269,11498,12132,13789,14149,
1085,1286,2630,3428,4056,5510,5991,6409,7720,8390,8543,11270,11499,12133,13790,14150,
1086,1287,2631,3429,4057,5511,5992,6410,7721,8391,8544,11271,11500,12134,13791,14151,
1087,1288,2632,3430,4058,5512,5993,6411,7722,8392,8545,11272,11501,12135,13792,14152,
1088,1289,2633,3431,4059,5513,5994,6412,7723,8393,8546,11273,11502,12136,13793,14153,
1089,1290,2634,3432,4060,5514,5995,6413,7724,8394,8547,11274,11503,12137,13794,14154,
1090,1291,2635,3433,4061,5515,5996,6414,7725,8395,8548,11275,11504,12138,13795,14155,
1091,1292,2636,3434,4062,5516,5997,6415,7726,8396,8549,11276,11505,12139,13796,14156,
1092,1293,2637,3435,4063,5517,5998,6416,7727,8397,8550,11277,11506,12140,13797,14157,
1093,1294,2638,3436,4064,5518,5999,6417,7728,8398,8551,11278,11507,12141,13798,14158,
1094,1295,2639,3437,4065,5519,6000,6418,7729,8399,8552,11279,11508,12142,13799,14159,
1095,1296,2640,3438,4066,5520,6001,6419,7730,8400,8553,11280,11509,12143,13800,14160,
1096,1297,2641,3439,4067,5521,6002,6420,7731,8401,8554,11281,11510,12144,13801,14161,
1097,1298,2642,3440,4068,5522,6003,6421,7732,8402,8555,11282,11511,12145,13802,14162,
1098,1299,2643,3441,4069,5523,6004,6422,7733,8403,8556,11283,11512,12146,13803,14163,
1099,1300,2644,3442,4070,5524,6005,6423,7734,8404,8557,11284,11513,12147,13804,14164,
1100,1301,2645,3443,4071,5525,6006,6424,7735,8405,8558,11285,11514,12148,13805,14165,
1101,1302,2646,3444,4072,5526,6007,6425,7736,8406,8559,11286,11515,12149,13806,14166,
1102,1303,2647,3445,4073,5527,6008,6426,7737,8407,8560,11287,11516,12150,13807,14167,
1103,1304,2648,3446,4074,5528,6009,6427,7738,8408,8561,11288,11517,12151,13808,14168,
1104,1305,2649,3447,4075,5529,6010,6428,7739,8409,8562,11289,11518,12152,13809,14169,
1105,1306,2650,3448,4076,5530,6011,6429,7740,8410,8563,11290,11519,12153,13810,14170,
1106,1307,2651,3449,4077,5531,6012,6430,7741,8411,8564,11160,11291,12154,13811,14171,
1107,1308,2652,3450,4078,5532,6013,6431,7742,8412,8565,11161,11292,12155,13812,14172,
1108,1309,2653,3451,4079,5533,6014,6432,7743,8413,8566,11162,11293,12156,13813,14173,
1109,1310,2654,3452,4080,5534,6015,6433,7744,8414,8567,11163,11294,12157,13814,14174,
1110,1311,2655,3453,4081,5535,6016,6434,7745,8415,8568,11164,11295,12158,13815,14175,
1111,1312,2656,3454,4082,5536,6017,6435,7746,8416,8569,11165,11296,12159,13816,14176,
1112,1313,2657,3455,4083,5537,6018,6436,7747,8417,8570,11166,11297,12160,13817,14177,
1113,1314,2658,3456,4084,5538,6019,6437,7748,8418,8571,11167,11298,12161,13818,14178,
1114,1315,2659,3457,4085,5539,6020,6438,7749,8419,8572,11168,11299,12162,13819,14179,
1115,1316,2660,3458,4086,5540,6021,6439,7750,8420,8573,11169,11300,12163,13820,14180,
1116,1317,2661,3459,4087,5541,6022,6440,7751,8421,8574,11170,11301,12164,13821,14181,
1117,1318,2662,3460,4088,5542,6023,6441,7752,8422,8575,11171,11302,12165,13822,14182,
1118,1319,2663,3461,4089,5543,6024,6442,7753,8423,8576,11172,11303,12166,13823,14183,
1119,1320,2664,3462,4090,5544,6025,6443,7754,8424,8577,11173,11304,12167,13824,14184,
1120,1321,2665,3463,4091,5545,6026,6444,7755,8425,8578,11174,11305,12168,13825,14185,
1121,1322,2666,3464,4092,5546,6027,6445,7756,8426,8579,11175,11306,12169,13826,14186,
1122,1323,2667,3465,4093,5547,6028,6446,7757,8427,8580,11176,11307,12170,13827,14187,
1123,1324,2668,3466,4094,5548,6029,6447,7758,8428,8581,11177,11308,12171,13828,14188,
1124,1325,2669,3467,4095,5549,6030,6448,7759,8429,8582,11178,11309,12172,13829,14189,
1125,1326,2670,3468,4096,5550,6031,6449,7760,8430,8583,11179,11310,12173,13830,14190,
1126,1327,2671,3469,4097,5551,6032,6450,7761,8431,8584,11180,11311,12174,13831,14191,
1127,1328,2672,3470,4098,5552,6033,6451,7762,8432,8585,11181,11312,12175,13832,14192,
1128,1329,2673,3471,4099,5553,6034,6452,7763,8433,8586,11182,11313,12176,13833,14193,
1129,1330,2674,3472,4100,5554,6035,6453,7764,8434,8587,11183,11314,12177,13834,14194,
1130,1331,2675,3473,4101,5555,6036,6454,7765,8435,8588,11184,11315,12178,13835,14195,
1131,1332,2676,3474,4102,5556,6037,6455,7766,8436,8589,11185,11316,12179,13836,14196,
1132,1333,2677,3475,4103,5557,6038,6456,7767,8437,8590,11186,11317,12180,13837,14197,
1133,1334,2678,3476,4104,5558,6039,6457,7768,8438,8591,11187,11318,12181,13838,14198,
1134,1335,2679,3477,4105,5559,6040,6458,7769,8439,8592,11188,11319,12182,13839,14199,
1135,1336,2680,3478,4106,5560,6041,6459,7770,8440,8593,11189,11320,12183,13840,14200,
1136,1337,2681,3479,4107,5561,6042,6460,7771,8441,8594,11190,11321,12184,13841,14201,
1137,1338,2682,3480,4108,5562,6043,6461,7772,8442,8595,11191,11322,12185,13842,14202,
1138,1339,2683,3481,4109,5563,6044,6462,7773,8443,8596,11192,11323,12186,13843,14203,
1139,1340,2684,3482,4110,5564,6045,6463,7774,8444,8597,11193,11324,12187,13844,14204,
1140,1341,2685,3483,4111,5565,6046,6464,7775,8445,8598,11194,11325,12188,13845,14205,
1141,1342,2686,3484,4112,5566,6047,6465,7776,8446,8599,11195,11326,12189,13846,14206,
1142,1343,2687,3485,4113,5567,6048,6466,7777,8447,8600,11196,11327,12190,13847,14207,
1143,1344,2688,3486,4114,5568,6049,6467,7778,8448,8601,11197,11328,12191,13848,14208,
1144,1345,2689,3487,4115,5569,6050,6468,7779,8449,8602,11198,11329,12192,13849,14209,
1145,1346,2690,3488,4116,5570,6051,6469,7780,8450,8603,11199,11330,12193,13850,14210,
1146,1347,2691,3489,4117,5571,6052,6470,7781,8451,8604,11200,11331,12194,13851,14211,
1147,1348,2692,3490,4118,5572,6053,6471,7782,8452,8605,11201,11332,12195,13852,14212,
1148,1349,2693,3491,4119,5573,6054,6472,7783,8453,8606,11202,11333,12196,13853,14213,
1149,1350,2694,3492,4120,5574,6055,6473,7784,8454,8607,11203,11334,12197,13854,14214,
1150,1351,2695,3493,4121,5575,6056,6474,7785,8455,8608,11204,11335,12198,13855,14215,
1151,1352,2696,3494,4122,5576,6057,6475,7786,8456,8609,11205,11336,12199,13856,14216,
1152,1353,2697,3495,4123,5577,6058,6476,7787,8457,8610,11206,11337,12200,13857,14217,
1153,1354,2698,3496,4124,5578,6059,6477,7788,8458,8611,11207,11338,12201,13858,14218,
1154,1355,2699,3497,4125,5579,6060,6478,7789,8459,8612,11208,11339,12202,13859,14219,
1155,1356,2700,3498,4126,5580,6061,6479,7790,8460,8613,11209,11340,12203,13860,14220,
1156,1357,2701,3499,4127,5581,6062,6120,7791,8461,8614,11210,11341,12204,13861,14221,
1157,1358,2702,3500,4128,5582,6063,6121,7792,8462,8615,11211,11342,12205,13862,14222,
1158,1359,2703,3501,4129,5583,6064,6122,7793,8463,8616,11212,11343,12206,13863,14223,
1159,1360,2704,3502,4130,5584,6065,6123,7794,8464,8617,11213,11344,12207,13864,14224,
1160,1361,2705,3503,4131,5585,6066,6124,7795,8465,8618,11214,11345,12208,13865,14225,
1161,1362,2706,3504,4132,5586,6067,6125,7796,8466,8619,11215,11346,12209,13866,14226,
1162,1363,2707,3505,4133,5587,6068,6126,7797,8467,8620,11216,11347,12210,13867,14227,
1163,1364,2708,3506,4134,5588,6069,6127,7798,8468,8621,11217,11348,12211,13868,14228,
1164,1365,2709,3507,4135,5589,6070,6128,7799,8469,8622,11218,11349,12212,13869,14229,
1165,1366,2710,3508,4136,5590,6071,6129,7800,8470,8623,11219,11350,12213,13870,14230,
1166,1367,2711,3509,4137,5591,6072,6130,7801,8471,8624,11220,11351,12214,13871,14231,
1167,1368,2712,3510,4138,5592,6073,6131,7802,8472,8625,11221,11352,12215,13872,14232,
1168,1369,2713,3511,4139,5593,6074,6132,7803,8473,8626,11222,11353,12216,13873,14233,
1169,1370,2714,3512,4140,5594,6075,6133,7804,8474,8627,11223,11354,12217,13874,14234,
1170,1371,2715,3513,4141,5595,6076,6134,7805,8475,8628,11224,11355,12218,13875,14235,
1171,1372,2716,3514,4142,5596,6077,6135,7806,8476,8629,11225,11356,12219,13876,14236,
1172,1373,2717,3515,4143,5597,6078,6136,7807,8477,8630,11226,11357,12220,13877,14237,
1173,1374,2718,3516,4144,5598,6079,6137,7808,8478,8631,11227,11358,12221,13878,14238,
1174,1375,2719,3517,4145,5599,6080,6138,7809,8479,8632,11228,11359,12222,13879,14239,
1175,1376,2720,3518,4146,5600,6081,6139,7810,8480,8633,11229,11360,12223,13880,14240,
1176,1377,2721,3519,4147,5601,6082,6140,7811,8481,8634,11230,11361,12224,13881,14241,
1177,1378,2722,3520,4148,5602,6083,6141,7812,8482,8635,11231,11362,12225,13882,14242,
1178,1379,2723,3521,4149,5603,6084,6142,7813,8483,8636,11232,11363,12226,13883,14243,
1179,1380,2724,3522,4150,5604,6085,6143,7814,8484,8637,11233,11364,12227,13884,14244,
1180,1381,2725,3523,4151,5605,6086,6144,7815,8485,8638,11234,11365,12228,13885,14245,
1181,1382,2726,3524,4152,5606,6087,6145,7816,8486,8639,11235,11366,12229,13886,14246,
1182,1383,2727,3525,4153,5607,6088,6146,7817,8280,8487,11236,11367,12230,13887,14247,
1183,1384,2728,3526,4154,5608,6089,6147,7818,8281,8488,11237,11368,12231,13888,14248,
1184,1385,2729,3527,4155,5609,6090,6148,7819,8282,8489,11238,11369,12232,13889,14249,
1185,1386,2730,3528,4156,5610,6091,6149,7820,8283,8490,11239,11370,12233,13890,14250,
1186,1387,2731,3529,4157,5611,6092,6150,7821,8284,8491,11240,11371,12234,13891,14251,
1187,1388,2732,3530,4158,5612,6093,6151,7822,8285,8492,11241,11372,12235,13892,14252,
1188,1389,2733,3531,4159,5613,6094,6152,7823,8286,8493,11242,11373,12236,13893,14253,
1189,1390,2734,3532,4160,5614,6095,6153,7824,8287,8494,11243,11374,12237,13894,14254,
1190,1391,2735,3533,4161,5615,6096,6154,7825,8288,8495,11244,11375,12238,13895,14255,
1191,1392,2736,3534,4162,5616,6097,6155,7826,8289,8496,11245,11376,12239,13896,14256,
1192,1393,2737,3535,4163,5617,6098,6156,7827,8290,8497,11246,11377,11880,13897,14257,
1193,1394,2738,3536,4164,5618,6099,6157,7828,8291,8498,11247,11378,11881,13898,14258,
1194,1395,2739,3537,4165,5619,6100,6158,7829,8292,8499,11248,11379,11882,13899,14259,
1195,1396,2740,3538,4166,5620,6101,6159,7830,8293,8500,11249,11380,11883,13900,14260,
1196,1397,2741,3539,4167,5621,6102,6160,7831,8294,8501,11250,11381,11884,13901,14261,
1197,1398,2742,3540,4168,5622,6103,6161,7832,8295,8502,11251,11382,11885,13902,14262,
1198,1399,2743,3541,4169,5623,6104,6162,7833,8296,8503,11252,11383,11886,13903,14263,
1199,1400,2744,3542,4170,5624,6105,6163,7834,8297,8504,11253,11384,11887,13904,14264,
1200,1401,2745,3543,4171,5625,6106,6164,7835,8298,8505,11254,11385,11888,13905,14265,
1201,1402,2746,3544,4172,5626,6107,6165,7836,8299,8506,11255,11386,11889,13906,14266,
1202,1403,2747,3545,4173,5627,6108,6166,7837,8300,8507,11256,11387,11890,13907,14267,
1203,1404,2748,3546,4174,5628,6109,6167,7838,8301,8508,11257,11388,11891,13908,14268,
1204,1405,2749,3547,4175,5629,6110,6168,7839,8302,8509,11258,11389,11892,13909,14269,
1205,1406,2750,3548,4176,5630,6111,6169,7840,8303,8510,11259,11390,11893,13910,14270,
1206,1407,2751,3549,4177,5631,6112,6170,7841,8304,8511,11260,11391,11894,13911,14271,
1207,1408,2752,3550,4178,5632,6113,6171,7842,8305,8512,11261,11392,11895,13912,14272,
1208,1409,2753,3551,4179,5633,6114,6172,7843,8306,8513,11262,11393,11896,13913,14273,
1209,1410,2754,3552,4180,5634,6115,6173,7844,8307,8514,11263,11394,11897,13914,14274,
1210,1411,2755,3553,4181,5635,6116,6174,7845,8308,8515,11264,11395,11898,13915,14275,
1211,1412,2756,3554,4182,5636,6117,6175,7846,8309,8516,11265,11396,11899,13916,14276,
1212,1413,2757,3555,4183,5637,6118,6176,7847,8310,8517,11266,11397,11900,13917,14277,
1213,1414,2758,3556,4184,5638,6119,6177,7848,8311,8518,11267,11398,11901,13918,14278,
1214,1415,2759,3557,4185,5639,5760,6178,7849,8312,8519,11268,11399,11902,13919,14279,
1215,1416,2760,3558,4186,5640,5761,6179,7850,8313,8520,11269,11400,11903,13920,14280,
1216,1417,2761,3559,4187,5641,5762,6180,7851,8314,8521,11270,11401,11904,13921,14281,
1217,1418,2762,3560,4188,5642,5763,6181,7852,8315,8522,11271,11402,11905,13922,14282,
1218,1419,2763,3561,4189,5643,5764,6182,7853,8316,8523,11272,11403,11906,13923,14283,
1219,1420,2764,3562,4190,5644,5765,6183,7854,8317,8524,11273,11404,11907,13924,14284,
1220,1421,2765,3563,4191,5645,5766,6184,7855,8318,8525,11274,11405,11908,13925,14285,
1221,1422,2766,3564,4192,5646,5767,6185,7856,8319,8526,11275,11406,11909,13926,14286,
1222,1423,2767,3565,4193,5647,5768,6186,7857,8320,8527,11276,11407,11910,13927,14287,
1223,1424,2768,3566,4194,5648,5769,6187,7858,8321,8528,11277,11408,11911,13928,14288,
1224,1425,2769,3567,4195,5649,5770,6188,7859,8322,8529,11278,11409,11912,13929,14289,
1225,1426,2770,3568,4196,5650,5771,6189,7860,8323,8530,11279,11410,11913,13930,14290,
1226,1427,2771,3569,4197,5651,5772,6190,7861,8324,8531,11280,11411,11914,13931,14291,
1227,1428,2772,3570,4198,5652,5773,6191,7862,8325,8532,11281,11412,11915,13932,14292,
1228,1429,2773,3571,4199,5653,5774,6192,7863,8326,8533,11282,11413,11916,13933,14293,
1229,1430,2774,3572,4200,5654,5775,6193,7864,8327,8534,11283,11414,11917,13934,14294,
1230,1431,2775,3573,4201,5655,5776,6194,7865,8328,8535,11284,11415,11918,13935,14295,
1231,1432,2776,3574,4202,5656,5777,6195,7866,8329,8536,11285,11416,11919,13936,14296,
1232,1433,2777,3575,4203,5657,5778,6196,7867,8330,8537,11286,11417,11920,13937,14297,
1233,1434,2778,3576,4204,5658,5779,6197,7868,8331,8538,11287,11418,11921,13938,14298,
1234,1435,2779,3577,4205,5659,5780,6198,7869,8332,8539,11288,11419,11922,13939,14299,
1235,1436,2780,3578,4206,5660,5781,6199,7870,8333,8540,11289,11420,11923,13940,14300,
1236,1437,2781,3579,4207,5661,5782,6200,7871,8334,8541,11290,11421,11924,13941,14301,
1237,1438,2782,3580,4208,5662,5783,6201,7872,8335,8542,11291,11422,11925,13942,14302,
1238,1439,2783,3581,4209,5663,5784,6202,7873,8336,8543,11292,11423,11926,13943,14303,
1080,1239,2784,3582,4210,5664,5785,6203,7874,8337,8544,11293,11424,11927,13944,14304,
1081,1240,2785,3583,4211,5665,5786,6204,7875,8338,8545,11294,11425,11928,13945,14305,
1082,1241,2786,3584,4212,5666,5787,6205,7876,8339,8546,11295,11426,11929,13946,14306,
1083,1242,2787,3585,4213,5667,5788,6206,7877,8340,8547,11296,11427,11930,13947,14307,
1084,1243,2788,3586,4214,5668,5789,6207,7878,8341,8548,11297,11428,11931,13948,14308,
1085,1244,2789,3587,4215,5669,5790,6208,7879,8342,8549,11298,11429,11932,13949,14309,
1086,1245,2790,3588,4216,5670,5791,6209,7880,8343,8550,11299,11430,11933,13950,14310,
1087,1246,2791,3589,4217,5671,5792,6210,7881,8344,8551,11300,11431,11934,13951,14311,
1088,1247,2792,3590,4218,5672,5793,6211,7882,8345,8552,11301,11432,11935,13952,14312,
1089,1248,2793,3591,4219,5673,5794,6212,7883,8346,8553,11302,11433,11936,13953,14313,
1090,1249,2794,3592,4220,5674,5795,6213,7884,8347,8554,11303,11434,11937,13954,14314,
1091,1250,2795,3593,4221,5675,5796,6214,7885,8348,8555,11304,11435,11938,13955,14315,
1092,1251,2796,3594,4222,5676,5797,6215,7886,8349,8556,11305,11436,11939,13956,14316,
1093,1252,2797,3595,4223,5677,5798,6216,7887,8350,8557,11306,11437,11940,13957,14317,
1094,1253,2798,3596,4224,5678,5799,6217,7888,8351,8558,11307,11438,11941,13958,14318,
1095,1254,2799,3597,4225,5679,5800,6218,7889,8352,8559,11308,11439,11942,13959,14319,
1096,1255,2800,3598,4226,5680,5801,6219,7890,8353,8560,11309,11440,11943,13960,14320,
1097,1256,2801,3599,4227,5681,5802,6220,7891,8354,8561,11310,11441,11944,13961,14321,
1098,1257,2802,3240,4228,5682,5803,6221,7892,8355,8562,11311,11442,11945,13962,14322,
1099,1258,2803,3241,4229,5683,5804,6222,7893,8356,8563,11312,11443,11946,13963,14323,
1100,1259,2804,3242,4230,5684,5805,6223,7894,8357,8564,11313,11444,11947,13964,14324,
1101,1260,2805,3243,4231,5685,5806,6224,7895,8358,8565,11314,11445,11948,13965,14325,
1102,1261,2806,3244,4232,5686,5807,6225,7896,8359,8566,11315,11446,11949,13966,14326,
1103,1262,2807,3245,4233,5687,5808,6226,7897,8360,8567,11316,11447,11950,13967,14327,
1104,1263,2808,3246,4234,5688,5809,6227,7898,8361,8568,11317,11448,11951,13968,14328,
1105,1264,2809,3247,4235,5689,5810,6228,7899,8362,8569,11318,11449,11952,13969,14329,
1106,1265,2810,3248,4236,5690,5811,6229,7900,8363,8570,11319,11450,11953,13970,14330,
1107,1266,2811,3249,4237,5691,5812,6230,7901,8364,8571,11320,11451,11954,13971,14331,
1108,1267,2812,3250,4238,5692,5813,6231,7902,8365,8572,11321,11452,11955,13972,14332,
1109,1268,2813,3251,4239,5693,5814,6232,7903,8366,8573,11322,11453,11956,13973,14333,
1110,1269,2814,3252,4240,5694,5815,6233,7904,8367,8574,11323,11454,11957,13974,14334,
1111,1270,2815,3253,4241,5695,5816,6234,7905,8368,8575,11324,11455,11958,13975,14335,
1112,1271,2816,3254,4242,5696,5817,6235,7906,8369,8576,11325,11456,11959,13976,14336,
1113,1272,2817,3255,4243,5697,5818,6236,7907,8370,8577,11326,11457,11960,13977,14337,
1114,1273,2818,3256,4244,5698,5819,6237,7908,8371,8578,11327,11458,11961,13978,14338,
1115,1274,2819,3257,4245,5699,5820,6238,7909,8372,8579,11328,11459,11962,13979,14339,
1116,1275,2820,3258,4246,5700,5821,6239,7910,8373,8580,11329,11460,11963,13980,14340,
1117,1276,2821,3259,4247,5701,5822,6240,7911,8374,8581,11330,11461,11964,13981,14341,
1118,1277,2822,3260,4248,5702,5823,6241,7912,8375,8582,11331,11462,11965,13982,14342,
1119,1278,2823,3261,4249,5703,5824,6242,7913,8376,8583,11332,11463,11966,13983,14343,
1120,1279,2824,3262,4250,5704,5825,6243,7914,8377,8584,11333,11464,11967,13984,14344,
1121,1280,2825,3263,4251,5705,5826,6244,7915,8378,8585,11334,11465,11968,13985,14345,
1122,1281,2826,3264,4252,5706,5827,6245,7916,8379,8586,11335,11466,11969,13986,14346,
1123,1282,2827,3265,4253,5707,5828,6246,7917,8380,8587,11336,11467,11970,13987,14347,
1124,1283,2828,3266,4254,5708,5829,6247,7918,8381,8588,11337,11468,11971,13988,14348,
1125,1284,2829,3267,4255,5709,5830,6248,7919,8382,8589,11338,11469,11972,13989,14349,
1126,1285,2830,3268,4256,5710,5831,6249,7560,8383,8590,11339,11470,11973,13990,14350,
1127,1286,2831,3269,4257,5711,5832,6250,7561,8384,8591,11340,11471,11974,13991,14351,
1128,1287,2832,3270,4258,5712,5833,6251,7562,8385,8592,11341,11472,11975,13992,14352,
1129,1288,2833,3271,4259,5713,5834,6252,7563,8386,8593,11342,11473,11976,13993,14353,
1130,1289,2834,3272,4260,5714,5835,6253,7564,8387,8594,11343,11474,11977,13994,14354,
1131,1290,2835,3273,4261,5715,5836,6254,7565,8388,8595,11344,11475,11978,13995,14355,
1132,1291,2836,3274,4262,5716,5837,6255,7566,8389,8596,11345,11476,11979,13996,14356,
1133,1292,2837,3275,4263,5717,5838,6256,7567,8390,8597,11346,11477,11980,13997,14357,
1134,1293,2838,3276,4264,5718,5839,6257,7568,8391,8598,11347,11478,11981,13998,14358,
1135,1294,2839,3277,4265,5719,5840,6258,7569,8392,8599,11348,11479,11982,13999,14359,
1136,1295,2840,3278,4266,5720,5841,6259,7570,8393,8600,11349,11480,11983,14000,14360,
1137,1296,2841,3279,4267,5721,5842,6260,7571,8394,8601,11350,11481,11984,14001,14361,
1138,1297,2842,3280,4268,5722,5843,6261,7572,8395,8602,11351,11482,11985,14002,14362,
1139,1298,2843,3281,4269,5723,5844,6262,7573,8396,8603,11352,11483,11986,14003,14363,
1140,1299,2844,3282,4270,5724,5845,6263,7574,8397,8604,11353,11484,11987,14004,14364,
1141,1300,2845,3283,4271,5725,5846,6264,7575,8398,8605,11354,11485,11988,14005,14365,
1142,1301,2846,3284,4272,5726,5847,6265,7576,8399,8606,11355,11486,11989,14006,14366,
1143,1302,2847,3285,4273,5727,5848,6266,7577,8400,8607,11356,11487,11990,14007,14367,
1144,1303,2848,3286,4274,5728,5849,6267,7578,8401,8608,11357,11488,11991,14008,14368,
1145,1304,2849,3287,4275,5729,5850,6268,7579,8402,8609,11358,11489,11992,14009,14369,
1146,1305,2850,3288,4276,5730,5851,6269,7580,8403,8610,11359,11490,11993,14010,14370,
1147,1306,2851,3289,4277,5731,5852,6270,7581,8404,8611,11360,11491,11994,14011,14371,
1148,1307,2852,3290,4278,5732,5853,6271,7582,8405,8612,11361,11492,11995,14012,14372,
1149,1308,2853,3291,4279,5733,5854,6272,7583,8406,8613,11362,11493,11996,14013,14373,
1150,1309,2854,3292,4280,5734,5855,6273,7584,8407,8614,11363,11494,11997,14014,14374,
1151,1310,2855,3293,4281,5735,5856,6274,7585,8408,8615,11364,11495,11998,14015,14375,
1152,1311,2856,3294,4282,5736,5857,6275,7586,8409,8616,11365,11496,11999,14016,14376,
1153,1312,2857,3295,4283,5737,5858,6276,7587,8410,8617,11366,11497,12000,14017,14377,
1154,1313,2858,3296,4284,5738,5859,6277,7588,8411,8618,11367,11498,12001,14018,14378,
1155,1314,2859,3297,4285,5739,5860,6278,7589,8412,8619,11368,11499,12002,14019,14379,
1156,1315,2860,3298,4286,5740,5861,6279,7590,8413,8620,11369,11500,12003,14020,14380,
1157,1316,2861,3299,4287,5741,5862,6280,7591,8414,8621,11370,11501,12004,14021,14381,
1158,1317,2862,3300,4288,5742,5863,6281,7592,8415,8622,11371,11502,12005,14022,14382,
1159,1318,2863,3301,4289,5743,5864,6282,7593,8416,8623,11372,11503,12006,14023,14383,
1160,1319,2864,3302,4290,5744,5865,6283,7594,8417,8624,11373,11504,12007,14024,14384,
1161,1320,2865,3303,4291,5745,5866,6284,7595,8418,8625,11374,11505,12008,14025,14385,
1162,1321,2866,3304,4292,5746,5867,6285,7596,8419,8626,11375,11506,12009,14026,14386,
1163,1322,2867,3305,4293,5747,5868,6286,7597,8420,8627,11376,11507,12010,14027,14387,
1164,1323,2868,3306,4294,5748,5869,6287,7598,8421,8628,11377,11508,12011,14028,14388,
1165,1324,2869,3307,4295,5749,5870,6288,7599,8422,8629,11378,11509,12012,14029,14389,
1166,1325,2870,3308,4296,5750,5871,6289,7600,8423,8630,11379,11510,12013,14030,14390,
1167,1326,2871,3309,4297,5751,5872,6290,7601,8424,8631,11380,11511,12014,14031,14391,
1168,1327,2872,3310,4298,5752,5873,6291,7602,8425,8632,11381,11512,12015,14032,14392,
1169,1328,2873,3311,4299,5753,5874,6292,7603,8426,8633,11382,11513,12016,14033,14393,
1170,1329,2874,3312,4300,5754,5875,6293,7604,8427,8634,11383,11514,12017,14034,14394,
1171,1330,2875,3313,4301,5755,5876,6294,7605,8428,8635,11384,11515,12018,14035,14395,
1172,1331,2876,3314,4302,5756,5877,6295,7606,8429,8636,11385,11516,12019,14036,14396,
1173,1332,2877,3315,4303,5757,5878,6296,7607,8430,8637,11386,11517,12020,14037,14397,
1174,1333,2878,3316,4304,5758,5879,6297,7608,8431,8638,11387,11518,12021,14038,14398,
1175,1334,2879,3317,4305,5759,5880,6298,7609,8432,8639,11388,11519,12022,14039,14399,
0,298,2778,2880,4400,5760,6829,7363,8640,9386,10026,11100,11520,12940,14040,14400,
1,299,2779,2881,4401,5761,6830,7364,8641,9387,10027,11101,11521,12941,14041,14401,
2,300,2780,2882,4402,5762,6831,7365,8642,9388,10028,11102,11522,12942,14042,14402,
3,301,2781,2883,4403,5763,6832,7366,8643,9389,10029,11103,11523,12943,14043,14403,
4,302,2782,2884,4404,5764,6833,7367,8644,9390,10030,11104,11524,12944,14044,14404,
5,303,2783,2885,4405,5765,6834,7368,8645,9391,10031,11105,11525,12945,14045,14405,
6,304,2784,2886,4406,5766,6835,7369,8646,9392,10032,11106,11526,12946,14046,14406,
7,305,2785,2887,4407,5767,6836,7370,8647,9393,10033,11107,11527,12947,14047,14407,
8,306,2786,2888,4408,5768,6837,7371,8648,9394,10034,11108,11528,12948,14048,14408,
9,307,2787,2889,4409,5769,6838,7372,8649,9395,10035,11109,11529,12949,14049,14409,
10,308,2788,2890,4410,5770,6839,7373,8650,9396,10036,11110,11530,12950,14050,14410,
11,309,2789,2891,4411,5771,6480,7374,8651,9397,10037,11111,11531,12951,14051,14411,
12,310,2790,2892,4412,5772,6481,7375,8652,9398,10038,11112,11532,12952,14052,14412,
13,311,2791,2893,4413,5773,6482,7376,8653,9399,10039,11113,11533,12953,14053,14413,
14,312,2792,2894,4414,5774,6483,7377,8654,9400,10040,11114,11534,12954,14054,14414,
15,313,2793,2895,4415,5775,6484,7378,8655,9401,10041,11115,11535,12955,14055,14415,
16,314,2794,2896,4416,5776,6485,7379,8656,9402,10042,11116,11536,12956,14056,14416,
17,315,2795,2897,4417,5777,6486,7380,8657,9403,10043,11117,11537,12957,14057,14417,
18,316,2796,2898,4418,5778,6487,7381,8658,9404,10044,11118,11538,12958,14058,14418,
19,317,2797,2899,4419,5779,6488,7382,8659,9405,10045,11119,11539,12959,14059,14419,
20,318,2798,2900,4420,5780,6489,7383,8660,9406,10046,11120,11540,12600,14060,14420,
21,319,2799,2901,4421,5781,6490,7384,8661,9407,10047,11121,11541,12601,14061,14421,
22,320,2800,2902,4422,5782,6491,7385,8662,9408,10048,11122,11542,12602,14062,14422,
23,321,2801,2903,4423,5783,6492,7386,8663,9409,10049,11123,11543,12603,14063,14423,
24,322,2802,2904,4424,5784,6493,7387,8664,9410,10050,11124,11544,12604,14064,14424,
25,323,2803,2905,4425,5785,6494,7388,8665,9411,10051,11125,11545,12605,14065,14425,
26,324,2804,2906,4426,5786,6495,7389,8666,9412,10052,11126,11546,12606,14066,14426,
27,325,2805,2907,4427,5787,6496,7390,8667,9413,10053,11127,11547,12607,14067,14427,
28,326,2806,2908,4428,5788,6497,7391,8668,9414,10054,11128,11548,12608,14068,14428,
29,327,2807,2909,4429,5789,6498,7392,8669,9415,10055,11129,11549,12609,14069,14429,
30,328,2808,2910,4430,5790,6499,7393,8670,9416,10056,11130,11550,12610,14070,14430,
31,329,2809,2911,4431,5791,6500,7394,8671,9417,10057,11131,11551,12611,14071,14431,
32,330,2810,2912,4432,5792,6501,7395,8672,9418,10058,11132,11552,12612,14072,14432,
33,331,2811,2913,4433,5793,6502,7396,8673,9419,10059,11133,11553,12613,14073,14433,
34,332,2812,2914,4434,5794,6503,7397,8674,9420,10060,11134,11554,12614,14074,14434,
35,333,2813,2915,4435,5795,6504,7398,8675,9421,10061,11135,11555,12615,14075,14435,
36,334,2814,2916,4436,5796,6505,7399,8676,9422,10062,11136,11556,12616,14076,14436,
37,335,2815,2917,4437,5797,6506,7400,8677,9423,10063,11137,11557,12617,14077,14437,
38,336,2816,2918,4438,5798,6507,7401,8678,9424,10064,11138,11558,12618,14078,14438,
39,337,2817,2919,4439,5799,6508,7402,8679,9425,10065,11139,11559,12619,14079,14439,
40,338,2818,2920,4440,5800,6509,7403,8680,9426,10066,11140,11560,12620,14080,14440,
41,339,2819,2921,4441,5801,6510,7404,8681,9427,10067,11141,11561,12621,14081,14441,
42,340,2820,2922,4442,5802,6511,7405,8682,9428,10068,11142,11562,12622,14082,14442,
43,341,2821,2923,4443,5803,6512,7406,8683,9429,10069,11143,11563,12623,14083,14443,
44,342,2822,2924,4444,5804,6513,7407,8684,9430,10070,11144,11564,12624,14084,14444,
45,343,2823,2925,4445,5805,6514,7408,8685,9431,10071,11145,11565,12625,14085,14445,
46,344,2824,2926,4446,5806,6515,7409,8686,9432,10072,11146,11566,12626,14086,14446,
47,345,2825,2927,4447,5807,6516,7410,8687,9433,10073,11147,11567,12627,14087,14447,
48,346,2826,2928,4448,5808,6517,7411,8688,9434,10074,11148,11568,12628,14088,14448,
49,347,2827,2929,4449,5809,6518,7412,8689,9435,10075,11149,11569,12629,14089,14449,
50,348,2828,2930,4450,5810,6519,7413,8690,9436,10076,11150,11570,12630,14090,14450,
51,349,2829,2931,4451,5811,6520,7414,8691,9437,10077,11151,11571,12631,14091,14451,
52,350,2830,2932,4452,5812,6521,7415,8692,9438,10078,11152,11572,12632,14092,14452,
53,351,2831,2933,4453,5813,6522,7416,8693,9439,10079,11153,11573,12633,14093,14453,
54,352,2832,2934,4454,5814,6523,7417,8694,9440,9720,11154,11574,12634,14094,14454,
55,353,2833,2935,4455,5815,6524,7418,8695,9441,9721,11155,11575,12635,14095,14455,
56,354,2834,2936,4456,5816,6525,7419,8696,9442,9722,11156,11576,12636,14096,14456,
57,355,2835,2937,4457,5817,6526,7420,8697,9443,9723,11157,11577,12637,14097,14457,
58,356,2836,2938,4458,5818,6527,7421,8698,9444,9724,11158,11578,12638,14098,14458,
59,357,2837,2939,4459,5819,6528,7422,8699,9445,9725,11159,11579,12639,14099,14459,
60,358,2838,2940,4460,5820,6529,7423,8700,9446,9726,10800,11580,12640,14100,14460,
61,359,2839,2941,4461,5821,6530,7424,8701,9447,9727,10801,11581,12641,14101,14461,
0,62,2840,2942,4462,5822,6531,7425,8702,9448,9728,10802,11582,12642,14102,14462,
1,63,2841,2943,4463,5823,6532,7426,8703,9449,9729,10803,11583,12643,14103,14463,
2,64,2842,2944,4464,5824,6533,7427,8704,9450,9730,10804,11584,12644,14104,14464,
3,65,2843,2945,4465,5825,6534,7428,8705,9451,9731,10805,11585,12645,14105,14465,
4,66,2844,2946,4466,5826,6535,7429,8706,9452,9732,10806,11586,12646,14106,14466,
5,67,2845,2947,4467,5827,6536,7430,8707,9453,9733,10807,11587,12647,14107,14467,
6,68,2846,2948,4468,5828,6537,7431,8708,9454,9734,10808,11588,12648,14108,14468,
7,69,2847,2949,4469,5829,6538,7432,8709,9455,9735,10809,11589,12649,14109,14469,
8,70,2848,2950,4470,5830,6539,7433,8710,9456,9736,10810,11590,12650,14110,14470,
9,71,2849,2951,4471,5831,6540,7434,8711,9457,9737,10811,11591,12651,14111,14471,
10,72,2850,2952,4472,5832,6541,7435,8712,9458,9738,10812,11592,12652,14112,14472,
11,73,2851,2953,4473,5833,6542,7436,8713,9459,9739,10813,11593,12653,14113,14473,
12,74,2852,2954,4474,5834,6543,7437,8714,9460,9740,10814,11594,12654,14114,14474,
13,75,2853,2955,4475,5835,6544,7438,8715,9461,9741,10815,11595,12655,14115,14475,
14,76,2854,2956,4476,5836,6545,7439,8716,9462,9742,10816,11596,12656,14116,14476,
15,77,2855,2957,4477,5837,6546,7440,8717,9463,9743,10817,11597,12657,14117,14477,
16,78,2856,2958,4478,5838,6547,7441,8718,9464,9744,10818,11598,12658,14118,14478,
17,79,2857,2959,4479,5839,6548,7442,8719,9465,9745,10819,11599,12659,14119,14479,
18,80,2858,2960,4480,5840,6549,7443,8720,9466,9746,10820,11600,12660,14120,14480,
19,81,2859,2961,4481,5841,6550,7444,8721,9467,9747,10821,11601,12661,14121,14481,
20,82,2860,2962,4482,5842,6551,7445,8722,9468,9748,10822,11602,12662,14122,14482,
21,83,2861,2963,4483,5843,6552,7446,8723,9469,9749,10823,11603,12663,14123,14483,
22,84,2862,2964,4484,5844,6553,7447,8724,9470,9750,10824,11604,12664,14124,14484,
23,85,2863,2965,4485,5845,6554,7448,8725,9471,9751,10825,11605,12665,14125,14485,
24,86,2864,2966,4486,5846,6555,7449,8726,9472,9752,10826,11606,12666,14126,14486,
25,87,2865,2967,4487,5847,6556,7450,8727,9473,9753,10827,11607,12667,14127,14487,
26,88,2866,2968,4488,5848,6557,7451,8728,9474,9754,10828,11608,12668,14128,14488,
27,89,2867,2969,4489,5849,6558,7452,8729,9475,9755,10829,11609,12669,14129,14489,
28,90,2868,2970,4490,5850,6559,7453,8730,9476,9756,10830,11610,12670,14130,14490,
29,91,2869,2971,4491,5851,6560,7454,8731,9477,9757,10831,11611,12671,14131,14491,
30,92,2870,2972,4492,5852,6561,7455,8732,9478,9758,10832,11612,12672,14132,14492,
31,93,2871,2973,4493,5853,6562,7456,8733,9479,9759,10833,11613,12673,14133,14493,
32,94,2872,2974,4494,5854,6563,7457,8734,9480,9760,10834,11614,12674,14134,14494,
33,95,2873,2975,4495,5855,6564,7458,8735,9481,9761,10835,11615,12675,14135,14495,
34,96,2874,2976,4496,5856,6565,7459,8736,9482,9762,10836,11616,12676,14136,14496,
35,97,2875,2977,4497,5857,6566,7460,8737,9483,9763,10837,11617,12677,14137,14497,
36,98,2876,2978,4498,5858,6567,7461,8738,9484,9764,10838,11618,12678,14138,14498,
37,99,2877,2979,4499,5859,6568,7462,8739,9485,9765,10839,11619,12679,14139,14499,
38,100,2878,2980,4500,5860,6569,7463,8740,9486,9766,10840,11620,12680,14140,14500,
39,101,2879,2981,4501,5861,6570,7464,8741,9487,9767,10841,11621,12681,14141,14501,
40,102,2520,2982,4502,5862,6571,7465,8742,9488,9768,10842,11622,12682,14142,14502,
41,103,2521,2983,4503,5863,6572,7466,8743,9489,9769,10843,11623,12683,14143,14503,
42,104,2522,2984,4504,5864,6573,7467,8744,9490,9770,10844,11624,12684,14144,14504,
43,105,2523,2985,4505,5865,6574,7468,8745,9491,9771,10845,11625,12685,14145,14505,
44,106,2524,2986,4506,5866,6575,7469,8746,9492,9772,10846,11626,12686,14146,14506,
45,107,2525,2987,4507,5867,6576,7470,8747,9493,9773,10847,11627,12687,14147,14507,
46,108,2526,2988,4508,5868,6577,7471,8748,9494,9774,10848,11628,12688,14148,14508,
47,109,2527,2989,4509,5869,6578,7472,8749,9495,9775,10849,11629,12689,14149,14509,
48,110,2528,2990,4510,5870,6579,7473,8750,9496,9776,10850,11630,12690,14150,14510,
49,111,2529,2991,4511,5871,6580,7474,8751,9497,9777,10851,11631,12691,14151,14511,
50,112,2530,2992,4512,5872,6581,7475,8752,9498,9778,10852,11632,12692,14152,14512,
51,113,2531,2993,4513,5873,6582,7476,8753,9499,9779,10853,11633,12693,14153,14513,
52,114,2532,2994,4514,5874,6583,7477,8754,9500,9780,10854,11634,12694,14154,14514,
53,115,2533,2995,4515,5875,6584,7478,8755,9501,9781,10855,11635,12695,14155,14515,
54,116,2534,2996,4516,5876,6585,7479,8756,9502,9782,10856,11636,12696,14156,14516,
55,117,2535,2997,4517,5877,6586,7480,8757,9503,9783,10857,11637,12697,14157,14517,
56,118,2536,2998,4518,5878,6587,7481,8758,9504,9784,10858,11638,12698,14158,14518,
57,119,2537,2999,4519,5879,6588,7482,8759,9505,9785,10859,11639,12699,14159,14519,
58,120,2538,3000,4520,5880,6589,7483,8760,9506,9786,10860,11640,12700,14160,14520,
59,121,2539,3001,4521,5881,6590,7484,8761,9507,9787,10861,11641,12701,14161,14521,
60,122,2540,3002,4522,5882,6591,7485,8762,9508,9788,10862,11642,12702,14162,14522,
61,123,2541,3003,4523,5883,6592,7486,8763,9509,9789,10863,11643,12703,14163,14523,
62,124,2542,3004,4524,5884,6593,7487,8764,9510,9790,10864,11644,12704,14164,14524,
63,125,2543,3005,4525,5885,6594,7488,8765,9511,9791,10865,11645,12705,14165,14525,
64,126,2544,3006,4526,5886,6595,7489,8766,9512,9792,10866,11646,12706,14166,14526,
65,127,2545,3007,4527,5887,6596,7490,8767,9513,9793,10867,11647,12707,14167,14527,
66,128,2546,3008,4528,5888,6597,7491,8768,9514,9794,10868,11648,12708,14168,14528,
67,129,2547,3009,4529,5889,6598,7492,8769,9515,9795,10869,11649,12709,14169,14529,
68,130,2548,3010,4530,5890,6599,7493,8770,9516,9796,10870,11650,12710,14170,14530,
69,131,2549,3011,4531,5891,6600,7494,8771,9517,9797,10871,11651,12711,14171,14531,
70,132,2550,3012,4532,5892,6601,7495,8772,9518,9798,10872,11652,12712,14172,14532,
71,133,2551,3013,4533,5893,6602,7496,8773,9519,9799,10873,11653,12713,14173,14533,
72,134,2552,3014,4534,5894,6603,7497,8774,9520,9800,10874,11654,12714,14174,14534,
73,135,2553,3015,4535,5895,6604,7498,8775,9521,9801,10875,11655,12715,14175,14535,
74,136,2554,3016,4536,5896,6605,7499,8776,9522,9802,10876,11656,12716,14176,14536,
75,137,2555,3017,4537,5897,6606,7500,8777,9523,9803,10877,11657,12717,14177,14537,
76,138,2556,3018,4538,5898,6607,7501,8778,9524,9804,10878,11658,12718,14178,14538,
77,139,2557,3019,4539,5899,6608,7502,8779,9525,9805,10879,11659,12719,14179,14539,
78,140,2558,3020,4540,5900,6609,7503,8780,9526,9806,10880,11660,12720,14180,14540,
79,141,2559,3021,4541,5901,6610,7504,8781,9527,9807,10881,11661,12721,14181,14541,
80,142,2560,3022,4542,5902,6611,7505,8782,9528,9808,10882,11662,12722,14182,14542,
81,143,2561,3023,4543,5903,6612,7506,8783,9529,9809,10883,11663,12723,14183,14543,
82,144,2562,3024,4544,5904,6613,7507,8784,9530,9810,10884,11664,12724,14184,14544,
83,145,2563,3025,4545,5905,6614,7508,8785,9531,9811,10885,11665,12725,14185,14545,
84,146,2564,3026,4546,5906,6615,7509,8786,9532,9812,10886,11666,12726,14186,14546,
85,147,2565,3027,4547,5907,6616,7510,8787,9533,9813,10887,11667,12727,14187,14547,
86,148,2566,3028,4548,5908,6617,7511,8788,9534,9814,10888,11668,12728,14188,14548,
87,149,2567,3029,4549,5909,6618,7512,8789,9535,9815,10889,11669,12729,14189,14549,
88,150,2568,3030,4550,5910,6619,7513,8790,9536,9816,10890,11670,12730,14190,14550,
89,151,2569,3031,4551,5911,6620,7514,8791,9537,9817,10891,11671,12731,14191,14551,
90,152,2570,3032,4552,5912,6621,7515,8792,9538,9818,10892,11672,12732,14192,14552,
91,153,2571,3033,4553,5913,6622,7516,8793,9539,9819,10893,11673,12733,14193,14553,
92,154,2572,3034,4554,5914,6623,7517,8794,9540,9820,10894,11674,12734,14194,14554,
93,155,2573,3035,4555,5915,6624,7518,8795,9541,9821,10895,11675,12735,14195,14555,
94,156,2574,3036,4556,5916,6625,7519,8796,9542,9822,10896,11676,12736,14196,14556,
95,157,2575,3037,4557,5917,6626,7520,8797,9543,9823,10897,11677,12737,14197,14557,
96,158,2576,3038,4558,5918,6627,7521,8798,9544,9824,10898,11678,12738,14198,14558,
97,159,2577,3039,4559,5919,6628,7522,8799,9545,9825,10899,11679,12739,14199,14559,
98,160,2578,3040,4560,5920,6629,7523,8800,9546,9826,10900,11680,12740,14200,14560,
99,161,2579,3041,4561,5921,6630,7524,8801,9547,9827,10901,11681,12741,14201,14561,
100,162,2580,3042,4562,5922,6631,7525,8802,9548,9828,10902,11682,12742,14202,14562,
101,163,2581,3043,4563,5923,6632,7526,8803,9549,9829,10903,11683,12743,14203,14563,
102,164,2582,3044,4564,5924,6633,7527,8804,9550,9830,10904,11684,12744,14204,14564,
103,165,2583,3045,4565,5925,6634,7528,8805,9551,9831,10905,11685,12745,14205,14565,
104,166,2584,3046,4566,5926,6635,7529,8806,9552,9832,10906,11686,12746,14206,14566,
105,167,2585,3047,4567,5927,6636,7530,8807,9553,9833,10907,11687,12747,14207,14567,
106,168,2586,3048,4568,5928,6637,7531,8808,9554,9834,10908,11688,12748,14208,14568,
107,169,2587,3049,4569,5929,6638,7532,8809,9555,9835,10909,11689,12749,14209,14569,
108,170,2588,3050,4570,5930,6639,7533,8810,9556,9836,10910,11690,12750,14210,14570,
109,171,2589,3051,4571,5931,6640,7534,8811,9557,9837,10911,11691,12751,14211,14571,
110,172,2590,3052,4572,5932,6641,7535,8812,9558,9838,10912,11692,12752,14212,14572,
111,173,2591,3053,4573,5933,6642,7536,8813,9559,9839,10913,11693,12753,14213,14573,
112,174,2592,3054,4574,5934,6643,7537,8814,9560,9840,10914,11694,12754,14214,14574,
113,175,2593,3055,4575,5935,6644,7538,8815,9561,9841,10915,11695,12755,14215,14575,
114,176,2594,3056,4576,5936,6645,7539,8816,9562,9842,10916,11696,12756,14216,14576,
115,177,2595,3057,4577,5937,6646,7540,8817,9563,9843,10917,11697,12757,14217,14577,
116,178,2596,3058,4578,5938,6647,7541,8818,9564,9844,10918,11698,12758,14218,14578,
117,179,2597,3059,4579,5939,6648,7542,8819,9565,9845,10919,11699,12759,14219,14579,
118,180,2598,3060,4580,5940,6649,7543,8820,9566,9846,10920,11700,12760,14220,14580,
119,181,2599,3061,4581,5941,6650,7544,8821,9567,9847,10921,11701,12761,14221,14581,
120,182,2600,3062,4582,5942,6651,7545,8822,9568,9848,10922,11702,12762,14222,14582,
121,183,2601,3063,4583,5943,6652,7546,8823,9569,9849,10923,11703,12763,14223,14583,
122,184,2602,3064,4584,5944,6653,7547,8824,9570,9850,10924,11704,12764,14224,14584,
123,185,2603,3065,4585,5945,6654,7548,8825,9571,9851,10925,11705,12765,14225,14585,
124,186,2604,3066,4586,5946,6655,7549,8826,9572,9852,10926,11706,12766,14226,14586,
125,187,2605,3067,4587,5947,6656,7550,8827,9573,9853,10927,11707,12767,14227,14587,
126,188,2606,3068,4588,5948,6657,7551,8828,9574,9854,10928,11708,12768,14228,14588,
127,189,2607,3069,4589,5949,6658,7552,8829,9575,9855,10929,11709,12769,14229,14589,
128,190,2608,3070,4590,5950,6659,7553,8830,9576,9856,10930,11710,12770,14230,14590,
129,191,2609,3071,4591,5951,6660,7554,8831,9577,9857,10931,11711,12771,14231,14591,
130,192,2610,3072,4592,5952,6661,7555,8832,9578,9858,10932,11712,12772,14232,14592,
131,193,2611,3073,4593,5953,6662,7556,8833,9579,9859,10933,11713,12773,14233,14593,
132,194,2612,3074,4594,5954,6663,7557,8834,9580,9860,10934,11714,12774,14234,14594,
133,195,2613,3075,4595,5955,6664,7558,8835,9581,9861,10935,11715,12775,14235,14595,
134,196,2614,3076,4596,5956,6665,7559,8836,9582,9862,10936,11716,12776,14236,14596,
135,197,2615,3077,4597,5957,6666,7200,8837,9583,9863,10937,11717,12777,14237,14597,
136,198,2616,3078,4598,5958,6667,7201,8838,9584,9864,10938,11718,12778,14238,14598,
137,199,2617,3079,4599,5959,6668,7202,8839,9585,9865,10939,11719,12779,14239,14599,
138,200,2618,3080,4600,5960,6669,7203,8840,9586,9866,10940,11720,12780,14240,14600,
139,201,2619,3081,4601,5961,6670,7204,8841,9587,9867,10941,11721,12781,14241,14601,
140,202,2620,3082,4602,5962,6671,7205,8842,9588,9868,10942,11722,12782,14242,14602,
141,203,2621,3083,4603,5963,6672,7206,8843,9589,9869,10943,11723,12783,14243,14603,
142,204,2622,3084,4604,5964,6673,7207,8844,9590,9870,10944,11724,12784,14244,14604,
143,205,2623,3085,4605,5965,6674,7208,8845,9591,9871,10945,11725,12785,14245,14605,
144,206,2624,3086,4606,5966,6675,7209,8846,9592,9872,10946,11726,12786,14246,14606,
145,207,2625,3087,4607,5967,6676,7210,8847,9593,9873,10947,11727,12787,14247,14607,
146,208,2626,3088,4608,5968,6677,7211,8848,9594,9874,10948,11728,12788,14248,14608,
147,209,2627,3089,4609,5969,6678,7212,8849,9595,9875,10949,11729,12789,14249,14609,
148,210,2628,3090,4610,5970,6679,7213,8850,9596,9876,10950,11730,12790,14250,14610,
149,211,2629,3091,4611,5971,6680,7214,8851,9597,9877,10951,11731,12791,14251,14611,
150,212,2630,3092,4612,5972,6681,7215,8852,9598,9878,10952,11732,12792,14252,14612,
151,213,2631,3093,4613,5973,6682,7216,8853,9599,9879,10953,11733,12793,14253,14613,
152,214,2632,3094,4614,5974,6683,7217,8854,9600,9880,10954,11734,12794,14254,14614,
153,215,2633,3095,4615,5975,6684,7218,8855,9601,9881,10955,11735,12795,14255,14615,
154,216,2634,3096,4616,5976,6685,7219,8856,9602,9882,10956,11736,12796,14256,14616,
155,217,2635,3097,4617,5977,6686,7220,8857,9603,9883,10957,11737,12797,14257,14617,
156,218,2636,3098,4618,5978,6687,7221,8858,9604,9884,10958,11738,12798,14258,14618,
157,219,2637,3099,4619,5979,6688,7222,8859,9605,9885,10959,11739,12799,14259,14619,
158,220,2638,3100,4620,5980,6689,7223,8860,9606,9886,10960,11740,12800,14260,14620,
159,221,2639,3101,4621,5981,6690,7224,8861,9607,9887,10961,11741,12801,14261,14621,
160,222,2640,3102,4622,5982,6691,7225,8862,9608,9888,10962,11742,12802,14262,14622,
161,223,2641,3103,4623,5983,6692,7226,8863,9609,9889,10963,11743,12803,14263,14623,
162,224,2642,3104,4624,5984,6693,7227,8864,9610,9890,10964,11744,12804,14264,14624,
163,225,2643,3105,4625,5985,6694,7228,8865,9611,9891,10965,11745,12805,14265,14625,
164,226,2644,3106,4626,5986,6695,7229,8866,9612,9892,10966,11746,12806,14266,14626,
165,227,2645,3107,4627,5987,6696,7230,8867,9613,9893,10967,11747,12807,14267,14627,
166,228,2646,3108,4628,5988,6697,7231,8868,9614,9894,10968,11748,12808,14268,14628,
167,229,2647,3109,4629,5989,6698,7232,8869,9615,9895,10969,11749,12809,14269,14629,
168,230,2648,3110,4630,5990,6699,7233,8870,9616,9896,10970,11750,12810,14270,14630,
169,231,2649,3111,4631,5991,6700,7234,8871,9617,9897,10971,11751,12811,14271,14631,
170,232,2650,3112,4632,5992,6701,7235,8872,9618,9898,10972,11752,12812,14272,14632,
171,233,2651,3113,4633,5993,6702,7236,8873,9619,9899,10973,11753,12813,14273,14633,
172,234,2652,3114,4634,5994,6703,7237,8874,9620,9900,10974,11754,12814,14274,14634,
173,235,2653,3115,4635,5995,6704,7238,8875,9621,9901,10975,11755,12815,14275,14635,
174,236,2654,3116,4636,5996,6705,7239,8876,9622,9902,10976,11756,12816,14276,14636,
175,237,2655,3117,4637,5997,6706,7240,8877,9623,9903,10977,11757,12817,14277,14637,
176,238,2656,3118,4638,5998,6707,7241,8878,9624,9904,10978,11758,12818,14278,14638,
177,239,2657,3119,4639,5999,6708,7242,8879,9625,9905,10979,11759,12819,14279,14639,
178,240,2658,3120,4640,6000,6709,7243,8880,9626,9906,10980,11760,12820,14280,14640,
179,241,2659,3121,4641,6001,6710,7244,8881,9627,9907,10981,11761,12821,14281,14641,
180,242,2660,3122,4642,6002,6711,7245,8882,9628,9908,10982,11762,12822,14282,14642,
181,243,2661,3123,4643,6003,6712,7246,8883,9629,9909,10983,11763,12823,14283,14643,
182,244,2662,3124,4644,6004,6713,7247,8884,9630,9910,10984,11764,12824,14284,14644,
183,245,2663,3125,4645,6005,6714,7248,8885,9631,9911,10985,11765,12825,14285,14645,
184,246,2664,3126,4646,6006,6715,7249,8886,9632,9912,10986,11766,12826,14286,14646,
185,247,2665,3127,4647,6007,6716,7250,8887,9633,9913,10987,11767,12827,14287,14647,
186,248,2666,3128,4648,6008,6717,7251,8888,9634,9914,10988,11768,12828,14288,14648,
187,249,2667,3129,4649,6009,6718,7252,8889,9635,9915,10989,11769,12829,14289,14649,
188,250,2668,3130,4650,6010,6719,7253,8890,9636,9916,10990,11770,12830,14290,14650,
189,251,2669,3131,4651,6011,6720,7254,8891,9637,9917,10991,11771,12831,14291,14651,
190,252,2670,3132,4652,6012,6721,7255,8892,9638,9918,10992,11772,12832,14292,14652,
191,253,2671,3133,4653,6013,6722,7256,8893,9639,9919,10993,11773,12833,14293,14653,
192,254,2672,3134,4654,6014,6723,7257,8894,9640,9920,10994,11774,12834,14294,14654,
193,255,2673,3135,4655,6015,6724,7258,8895,9641,9921,10995,11775,12835,14295,14655,
194,256,2674,3136,4656,6016,6725,7259,8896,9642,9922,10996,11776,12836,14296,14656,
195,257,2675,3137,4657,6017,6726,7260,8897,9643,9923,10997,11777,12837,14297,14657,
196,258,2676,3138,4658,6018,6727,7261,8898,9644,9924,10998,11778,12838,14298,14658,
197,259,2677,3139,4659,6019,6728,7262,8899,9645,9925,10999,11779,12839,14299,14659,
198,260,2678,3140,4660,6020,6729,7263,8900,9646,9926,11000,11780,12840,14300,14660,
199,261,2679,3141,4661,6021,6730,7264,8901,9647,9927,11001,11781,12841,14301,14661,
200,262,2680,3142,4662,6022,6731,7265,8902,9648,9928,11002,11782,12842,14302,14662,
201,263,2681,3143,4663,6023,6732,7266,8903,9649,9929,11003,11783,12843,14303,14663,
202,264,2682,3144,4664,6024,6733,7267,8904,9650,9930,11004,11784,12844,14304,14664,
203,265,2683,3145,4665,6025,6734,7268,8905,9651,9931,11005,11785,12845,14305,14665,
204,266,2684,3146,4666,6026,6735,7269,8906,9652,9932,11006,11786,12846,14306,14666,
205,267,2685,3147,4667,6027,6736,7270,8907,9653,9933,11007,11787,12847,14307,14667,
206,268,2686,3148,4668,6028,6737,7271,8908,9654,9934,11008,11788,12848,14308,14668,
207,269,2687,3149,4669,6029,6738,7272,8909,9655,9935,11009,11789,12849,14309,14669,
208,270,2688,3150,4670,6030,6739,7273,8910,9656,9936,11010,11790,12850,14310,14670,
209,271,2689,3151,4671,6031,6740,7274,8911,9657,9937,11011,11791,12851,14311,14671,
210,272,2690,3152,4672,6032,6741,7275,8912,9658,9938,11012,11792,12852,14312,14672,
211,273,2691,3153,4673,6033,6742,7276,8913,9659,9939,11013,11793,12853,14313,14673,
212,274,2692,3154,4674,6034,6743,7277,8914,9660,9940,11014,11794,12854,14314,14674,
213,275,2693,3155,4675,6035,6744,7278,8915,9661,9941,11015,11795,12855,14315,14675,
214,276,2694,3156,4676,6036,6745,7279,8916,9662,9942,11016,11796,12856,14316,14676,
215,277,2695,3157,4677,6037,6746,7280,8917,9663,9943,11017,11797,12857,14317,14677,
216,278,2696,3158,4678,6038,6747,7281,8918,9664,9944,11018,11798,12858,14318,14678,
217,279,2697,3159,4679,6039,6748,7282,8919,9665,9945,11019,11799,12859,14319,14679,
218,280,2698,3160,4320,6040,6749,7283,8920,9666,9946,11020,11800,12860,14320,14680,
219,281,2699,3161,4321,6041,6750,7284,8921,9667,9947,11021,11801,12861,14321,14681,
220,282,2700,3162,4322,6042,6751,7285,8922,9668,9948,11022,11802,12862,14322,14682,
221,283,2701,3163,4323,6043,6752,7286,8923,9669,9949,11023,11803,12863,14323,14683,
222,284,2702,3164,4324,6044,6753,7287,8924,9670,9950,11024,11804,12864,14324,14684,
223,285,2703,3165,4325,6045,6754,7288,8925,9671,9951,11025,11805,12865,14325,14685,
224,286,2704,3166,4326,6046,6755,7289,8926,9672,9952,11026,11806,12866,14326,14686,
225,287,2705,3167,4327,6047,6756,7290,8927,9673,9953,11027,11807,12867,14327,14687,
226,288,2706,3168,4328,6048,6757,7291,8928,9674,9954,11028,11808,12868,14328,14688,
227,289,2707,3169,4329,6049,6758,7292,8929,9675,9955,11029,11809,12869,14329,14689,
228,290,2708,3170,4330,6050,6759,7293,8930,9676,9956,11030,11810,12870,14330,14690,
229,291,2709,3171,4331,6051,6760,7294,8931,9677,9957,11031,11811,12871,14331,14691,
230,292,2710,3172,4332,6052,6761,7295,8932,9678,9958,11032,11812,12872,14332,14692,
231,293,2711,3173,4333,6053,6762,7296,8933,9679,9959,11033,11813,12873,14333,14693,
232,294,2712,3174,4334,6054,6763,7297,8934,9680,9960,11034,11814,12874,14334,14694,
233,295,2713,3175,4335,6055,6764,7298,8935,9681,9961,11035,11815,12875,14335,14695,
234,296,2714,3176,4336,6056,6765,7299,8936,9682,9962,11036,11816,12876,14336,14696,
235,297,2715,3177,4337,6057,6766,7300,8937,9683,9963,11037,11817,12877,14337,14697,
236,298,2716,3178,4338,6058,6767,7301,8938,9684,9964,11038,11818,12878,14338,14698,
237,299,2717,3179,4339,6059,6768,7302,8939,9685,9965,11039,11819,12879,14339,14699,
238,300,2718,3180,4340,6060,6769,7303,8940,9686,9966,11040,11820,12880,14340,14700,
239,301,2719,3181,4341,6061,6770,7304,8941,9687,9967,11041,11821,12881,14341,14701,
240,302,2720,3182,4342,6062,6771,7305,8942,9688,9968,11042,11822,12882,14342,14702,
241,303,2721,3183,4343,6063,6772,7306,8943,9689,9969,11043,11823,12883,14343,14703,
242,304,2722,3184,4344,6064,6773,7307,8944,9690,9970,11044,11824,12884,14344,14704,
243,305,2723,3185,4345,6065,6774,7308,8945,9691,9971,11045,11825,12885,14345,14705,
244,306,2724,3186,4346,6066,6775,7309,8946,9692,9972,11046,11826,12886,14346,14706,
245,307,2725,3187,4347,6067,6776,7310,8947,9693,9973,11047,11827,12887,14347,14707,
246,308,2726,3188,4348,6068,6777,7311,8948,9694,9974,11048,11828,12888,14348,14708,
247,309,2727,3189,4349,6069,6778,7312,8949,9695,9975,11049,11829,12889,14349,14709,
248,310,2728,3190,4350,6070,6779,7313,8950,9696,9976,11050,11830,12890,14350,14710,
249,311,2729,3191,4351,6071,6780,7314,8951,9697,9977,11051,11831,12891,14351,14711,
250,312,2730,3192,4352,6072,6781,7315,8952,9698,9978,11052,11832,12892,14352,14712,
251,313,2731,3193,4353,6073,6782,7316,8953,9699,9979,11053,11833,12893,14353,14713,
252,314,2732,3194,4354,6074,6783,7317,8954,9700,9980,11054,11834,12894,14354,14714,
253,315,2733,3195,4355,6075,6784,7318,8955,9701,9981,11055,11835,12895,14355,14715,
254,316,2734,3196,4356,6076,6785,7319,8956,9702,9982,11056,11836,12896,14356,14716,
255,317,2735,3197,4357,6077,6786,7320,8957,9703,9983,11057,11837,12897,14357,14717,
256,318,2736,3198,4358,6078,6787,7321,8958,9704,9984,11058,11838,12898,14358,14718,
257,319,2737,3199,4359,6079,6788,7322,8959,9705,9985,11059,11839,12899,14359,14719,
258,320,2738,3200,4360,6080,6789,7323,8960,9706,9986,11060,11840,12900,14360,14720,
259,321,2739,3201,4361,6081,6790,7324,8961,9707,9987,11061,11841,12901,14361,14721,
260,322,2740,3202,4362,6082,6791,7325,8962,9708,9988,11062,11842,12902,14362,14722,
261,323,2741,3203,4363,6083,6792,7326,8963,9709,9989,11063,11843,12903,14363,14723,
262,324,2742,3204,4364,6084,6793,7327,8964,9710,9990,11064,11844,12904,14364,14724,
263,325,2743,3205,4365,6085,6794,7328,8965,9711,9991,11065,11845,12905,14365,14725,
264,326,2744,3206,4366,6086,6795,7329,8966,9712,9992,11066,11846,12906,14366,14726,
265,327,2745,3207,4367,6087,6796,7330,8967,9713,9993,11067,11847,12907,14367,14727,
266,328,2746,3208,4368,6088,6797,7331,8968,9714,9994,11068,11848,12908,14368,14728,
267,329,2747,3209,4369,6089,6798,7332,8969,9715,9995,11069,11849,12909,14369,14729,
268,330,2748,3210,4370,6090,6799,7333,8970,9716,9996,11070,11850,12910,14370,14730,
269,331,2749,3211,4371,6091,6800,7334,8971,9717,9997,11071,11851,12911,14371,14731,
270,332,2750,3212,4372,6092,6801,7335,8972,9718,9998,11072,11852,12912,14372,14732,
271,333,2751,3213,4373,6093,6802,7336,8973,9719,9999,11073,11853,12913,14373,14733,
272,334,2752,3214,4374,6094,6803,7337,8974,9360,10000,11074,11854,12914,14374,14734,
273,335,2753,3215,4375,6095,6804,7338,8975,9361,10001,11075,11855,12915,14375,14735,
274,336,2754,3216,4376,6096,6805,7339,8976,9362,10002,11076,11856,12916,14376,14736,
275,337,2755,3217,4377,6097,6806,7340,8977,9363,10003,11077,11857,12917,14377,14737,
276,338,2756,3218,4378,6098,6807,7341,8978,9364,10004,11078,11858,12918,14378,14738,
277,339,2757,3219,4379,6099,6808,7342,8979,9365,10005,11079,11859,12919,14379,14739,
278,340,2758,3220,4380,6100,6809,7343,8980,9366,10006,11080,11860,12920,14380,14740,
279,341,2759,3221,4381,6101,6810,7344,8981,9367,10007,11081,11861,12921,14381,14741,
280,342,2760,3222,4382,6102,6811,7345,8982,9368,10008,11082,11862,12922,14382,14742,
281,343,2761,3223,4383,6103,6812,7346,8983,9369,10009,11083,11863,12923,14383,14743,
282,344,2762,3224,4384,6104,6813,7347,8984,9370,10010,11084,11864,12924,14384,14744,
283,345,2763,3225,4385,6105,6814,7348,8985,9371,10011,11085,11865,12925,14385,14745,
284,346,2764,3226,4386,6106,6815,7349,8986,9372,10012,11086,11866,12926,14386,14746,
285,347,2765,3227,4387,6107,6816,7350,8987,9373,10013,11087,11867,12927,14387,14747,
286,348,2766,3228,4388,6108,6817,7351,8988,9374,10014,11088,11868,12928,14388,14748,
287,349,2767,3229,4389,6109,6818,7352,8989,9375,10015,11089,11869,12929,14389,14749,
288,350,2768,3230,4390,6110,6819,7353,8990,9376,10016,11090,11870,12930,14390,14750,
289,351,2769,3231,4391,6111,6820,7354,8991,9377,10017,11091,11871,12931,14391,14751,
290,352,2770,3232,4392,6112,6821,7355,8992,9378,10018,11092,11872,12932,14392,14752,
291,353,2771,3233,4393,6113,6822,7356,8993,9379,10019,11093,11873,12933,14393,14753,
292,354,2772,3234,4394,6114,6823,7357,8994,9380,10020,11094,11874,12934,14394,14754,
293,355,2773,3235,4395,6115,6824,7358,8995,9381,10021,11095,11875,12935,14395,14755,
294,356,2774,3236,4396,6116,6825,7359,8996,9382,10022,11096,11876,12936,14396,14756,
295,357,2775,3237,4397,6117,6826,7360,8997,9383,10023,11097,11877,12937,14397,14757,
296,358,2776,3238,4398,6118,6827,7361,8998,9384,10024,11098,11878,12938,14398,14758,
297,359,2777,3239,4399,6119,6828,7362,8999,9385,10025,11099,11879,12939,14399,14759,
47,247,271,360,1774,2227,3240,3840,6120,6414,6922,9000,9238,10412,11880,12232,12990,14400,14760,
48,248,272,361,1775,2228,3241,3841,6121,6415,6923,9001,9239,10413,11881,12233,12991,14401,14761,
49,249,273,362,1776,2229,3242,3842,6122,6416,6924,9002,9240,10414,11882,12234,12992,14402,14762,
50,250,274,363,1777,2230,3243,3843,6123,6417,6925,9003,9241,10415,11883,12235,12993,14403,14763,
51,251,275,364,1778,2231,3244,3844,6124,6418,6926,9004,9242,10416,11884,12236,12994,14404,14764,
52,252,276,365,1779,2232,3245,3845,6125,6419,6927,9005,9243,10417,11885,12237,12995,14405,14765,
53,253,277,366,1780,2233,3246,3846,6126,6420,6928,9006,9244,10418,11886,12238,12996,14406,14766,
54,254,278,367,1781,2234,3247,3847,6127,6421,6929,9007,9245,10419,11887,12239,12997,14407,14767,
55,255,279,368,1782,2235,3248,3848,6128,6422,6930,9008,9246,10420,11880,11888,12998,14408,14768,
56,256,280,369,1783,2236,3249,3849,6129,6423,6931,9009,9247,10421,11881,11889,12999,14409,14769,
57,257,281,370,1784,2237,3250,3850,6130,6424,6932,9010,9248,10422,11882,11890,13000,14410,14770,
58,258,282,371,1785,2238,3251,3851,6131,6425,6933,9011,9249,10423,11883,11891,13001,14411,14771,
59,259,283,372,1786,2239,3252,3852,6132,6426,6934,9012,9250,10424,11884,11892,13002,14412,14772,
60,260,284,373,1787,2240,3253,3853,6133,6427,6935,9013,9251,10425,11885,11893,13003,14413,14773,
61,261,285,374,1788,2241,3254,3854,6134,6428,6936,9014,9252,10426,11886,11894,13004,14414,14774,
62,262,286,375,1789,2242,3255,3855,6135,6429,6937,9015,9253,10427,11887,11895,13005,14415,14775,
63,263,287,376,1790,2243,3256,3856,6136,6430,6938,9016,9254,10428,11888,11896,13006,14416,14776,
64,264,288,377,1791,2244,3257,3857,6137,6431,6939,9017,9255,10429,11889,11897,13007,14417,14777,
65,265,289,378,1792,2245,3258,3858,6138,6432,6940,9018,9256,10430,11890,11898,13008,14418,14778,
66,266,290,379,1793,2246,3259,3859,6139,6433,6941,9019,9257,10431,11891,11899,13009,14419,14779,
67,267,291,380,1794,2247,3260,3860,6140,6434,6942,9020,9258,10432,11892,11900,13010,14420,14780,
68,268,292,381,1795,2248,3261,3861,6141,6435,6943,9021,9259,10433,11893,11901,13011,14421,14781,
69,269,293,382,1796,2249,3262,3862,6142,6436,6944,9022,9260,10434,11894,11902,13012,14422,14782,
70,270,294,383,1797,2250,3263,3863,6143,6437,6945,9023,9261,10435,11895,11903,13013,14423,14783,
71,271,295,384,1798,2251,3264,3864,6144,6438,6946,9024,9262,10436,11896,11904,13014,14424,14784,
72,272,296,385,1799,2252,3265,3865,6145,6439,6947,9025,9263,10437,11897,11905,13015,14425,14785,
73,273,297,386,1440,2253,3266,3866,6146,6440,6948,9026,9264,10438,11898,11906,13016,14426,14786,
74,274,298,387,1441,2254,3267,3867,6147,6441,6949,9027,9265,10439,11899,11907,13017,14427,14787,
75,275,299,388,1442,2255,3268,3868,6148,6442,6950,9028,9266,10080,11900,11908,13018,14428,14788,
76,276,300,389,1443,2256,3269,3869,6149,6443,6951,9029,9267,10081,11901,11909,13019,14429,14789,
77,277,301,390,1444,2257,3270,3870,6150,6444,6952,9030,9268,10082,11902,11910,13020,14430,14790,
78,278,302,391,1445,2258,3271,3871,6151,6445,6953,9031,9269,10083,11903,11911,13021,14431,14791,
79,279,303,392,1446,2259,3272,3872,6152,6446,6954,9032,9270,10084,11904,11912,13022,14432,14792,
80,280,304,393,1447,2260,3273,3873,6153,6447,6955,9033,9271,10085,11905,11913,13023,14433,14793,
81,281,305,394,1448,2261,3274,3874,6154,6448,6956,9034,9272,10086,11906,11914,13024,14434,14794,
82,282,306,395,1449,2262,3275,3875,6155,6449,6957,9035,9273,10087,11907,11915,13025,14435,14795,
83,283,307,396,1450,2263,3276,3876,6156,6450,6958,9036,9274,10088,11908,11916,13026,14436,14796,
84,284,308,397,1451,2264,3277,3877,6157,6451,6959,9037,9275,10089,11909,11917,13027,14437,14797,
85,285,309,398,1452,2265,3278,3878,6158,6452,6960,9038,9276,10090,11910,11918,13028,14438,14798,
86,286,310,399,1453,2266,3279,3879,6159,6453,6961,9039,9277,10091,11911,11919,13029,14439,14799,
87,287,311,400,1454,2267,3280,3880,6160,6454,6962,9040,9278,10092,11912,11920,13030,14440,14800,
88,288,312,401,1455,2268,3281,3881,6161,6455,6963,9041,9279,10093,11913,11921,13031,14441,14801,
89,289,313,402,1456,2269,3282,3882,6162,6456,6964,9042,9280,10094,11914,11922,13032,14442,14802,
90,290,314,403,1457,2270,3283,3883,6163,6457,6965,9043,9281,10095,11915,11923,13033,14443,14803,
91,291,315,404,1458,2271,3284,3884,6164,6458,6966,9044,9282,10096,11916,11924,13034,14444,14804,
92,292,316,405,1459,2272,3285,3885,6165,6459,6967,9045,9283,10097,11917,11925,13035,14445,14805,
93,293,317,406,1460,2273,3286,3886,6166,6460,6968,9046,9284,10098,11918,11926,13036,14446,14806,
94,294,318,407,1461,2274,3287,3887,6167,6461,6969,9047,9285,10099,11919,11927,13037,14447,14807,
95,295,319,408,1462,2275,3288,3888,6168,6462,6970,9048,9286,10100,11920,11928,13038,14448,14808,
96,296,320,409,1463,2276,3289,3889,6169,6463,6971,9049,9287,10101,11921,11929,13039,14449,14809,
97,297,321,410,1464,2277,3290,3890,6170,6464,6972,9050,9288,10102,11922,11930,13040,14450,14810,
98,298,322,411,1465,2278,3291,3891,6171,6465,6973,9051,9289,10103,11923,11931,13041,14451,14811,
99,299,323,412,1466,2279,3292,3892,6172,6466,6974,9052,9290,10104,11924,11932,13042,14452,14812,
100,300,324,413,1467,2280,3293,3893,6173,6467,6975,9053,9291,10105,11925,11933,13043,14453,14813,
101,301,325,414,1468,2281,3294,3894,6174,6468,6976,9054,9292,10106,11926,11934,13044,14454,14814,
102,302,326,415,1469,2282,3295,3895,6175,6469,6977,9055,9293,10107,11927,11935,13045,14455,14815,
103,303,327,416,1470,2283,3296,3896,6176,6470,6978,9056,9294,10108,11928,11936,13046,14456,14816,
104,304,328,417,1471,2284,3297,3897,6177,6471,6979,9057,9295,10109,11929,11937,13047,14457,14817,
105,305,329,418,1472,2285,3298,3898,6178,6472,6980,9058,9296,10110,11930,11938,13048,14458,14818,
106,306,330,419,1473,2286,3299,3899,6179,6473,6981,9059,9297,10111,11931,11939,13049,14459,14819,
107,307,331,420,1474,2287,3300,3900,6180,6474,6982,9060,9298,10112,11932,11940,13050,14460,14820,
108,308,332,421,1475,2288,3301,3901,6181,6475,6983,9061,9299,10113,11933,11941,13051,14461,14821,
109,309,333,422,1476,2289,3302,3902,6182,6476,6984,9062,9300,10114,11934,11942,13052,14462,14822,
110,310,334,423,1477,2290,3303,3903,6183,6477,6985,9063,9301,10115,11935,11943,13053,14463,14823,
111,311,335,424,1478,2291,3304,3904,6184,6478,6986,9064,9302,10116,11936,11944,13054,14464,14824,
112,312,336,425,1479,2292,3305,3905,6185,6479,6987,9065,9303,10117,11937,11945,13055,14465,14825,
113,313,337,426,1480,2293,3306,3906,6120,6186,6988,9066,9304,10118,11938,11946,13056,14466,14826,
114,314,338,427,1481,2294,3307,3907,6121,6187,6989,9067,9305,10119,11939,11947,13057,14467,14827,
115,315,339,428,1482,2295,3308,3908,6122,6188,6990,9068,9306,10120,11940,11948,13058,14468,14828,
116,316,340,429,1483,2296,3309,3909,6123,6189,6991,9069,9307,10121,11941,11949,13059,14469,14829,
117,317,341,430,1484,2297,3310,3910,6124,6190,6992,9070,9308,10122,11942,11950,13060,14470,14830,
118,318,342,431,1485,2298,3311,3911,6125,6191,6993,9071,9309,10123,11943,11951,13061,14471,14831,
119,319,343,432,1486,2299,3312,3912,6126,6192,6994,9072,9310,10124,11944,11952,13062,14472,14832,
120,320,344,433,1487,2300,3313,3913,6127,6193,6995,9073,9311,10125,11945,11953,13063,14473,14833,
121,321,345,434,1488,2301,3314,3914,6128,6194,6996,9074,9312,10126,11946,11954,13064,14474,14834,
122,322,346,435,1489,2302,3315,3915,6129,6195,6997,9075,9313,10127,11947,11955,13065,14475,14835,
123,323,347,436,1490,2303,3316,3916,6130,6196,6998,9076,9314,10128,11948,11956,13066,14476,14836,
124,324,348,437,1491,2304,3317,3917,6131,6197,6999,9077,9315,10129,11949,11957,13067,14477,14837,
125,325,349,438,1492,2305,3318,3918,6132,6198,7000,9078,9316,10130,11950,11958,13068,14478,14838,
126,326,350,439,1493,2306,3319,3919,6133,6199,7001,9079,9317,10131,11951,11959,13069,14479,14839,
127,327,351,440,1494,2307,3320,3920,6134,6200,7002,9080,9318,10132,11952,11960,13070,14480,14840,
128,328,352,441,1495,2308,3321,3921,6135,6201,7003,9081,9319,10133,11953,11961,13071,14481,14841,
129,329,353,442,1496,2309,3322,3922,6136,6202,7004,9082,9320,10134,11954,11962,13072,14482,14842,
130,330,354,443,1497,2310,3323,3923,6137,6203,7005,9083,9321,10135,11955,11963,13073,14483,14843,
131,331,355,444,1498,2311,3324,3924,6138,6204,7006,9084,9322,10136,11956,11964,13074,14484,14844,
132,332,356,445,1499,2312,3325,3925,6139,6205,7007,9085,9323,10137,11957,11965,13075,14485,14845,
133,333,357,446,1500,2313,3326,3926,6140,6206,7008,9086,9324,10138,11958,11966,13076,14486,14846,
134,334,358,447,1501,2314,3327,3927,6141,6207,7009,9087,9325,10139,11959,11967,13077,14487,14847,
135,335,359,448,1502,2315,3328,3928,6142,6208,7010,9088,9326,10140,11960,11968,13078,14488,14848,
0,136,336,449,1503,2316,3329,3929,6143,6209,7011,9089,9327,10141,11961,11969,13079,14489,14849,
1,137,337,450,1504,2317,3330,3930,6144,6210,7012,9090,9328,10142,11962,11970,13080,14490,14850,
2,138,338,451,1505,2318,3331,3931,6145,6211,7013,9091,9329,10143,11963,11971,13081,14491,14851,
3,139,339,452,1506,2319,3332,3932,6146,6212,7014,9092,9330,10144,11964,11972,13082,14492,14852,
4,140,340,453,1507,2320,3333,3933,6147,6213,7015,9093,9331,10145,11965,11973,13083,14493,14853,
5,141,341,454,1508,2321,3334,3934,6148,6214,7016,9094,9332,10146,11966,11974,13084,14494,14854,
6,142,342,455,1509,2322,3335,3935,6149,6215,7017,9095,9333,10147,11967,11975,13085,14495,14855,
7,143,343,456,1510,2323,3336,3936,6150,6216,7018,9096,9334,10148,11968,11976,13086,14496,14856,
8,144,344,457,1511,2324,3337,3937,6151,6217,7019,9097,9335,10149,11969,11977,13087,14497,14857,
9,145,345,458,1512,2325,3338,3938,6152,6218,7020,9098,9336,10150,11970,11978,13088,14498,14858,
10,146,346,459,1513,2326,3339,3939,6153,6219,7021,9099,9337,10151,11971,11979,13089,14499,14859,
11,147,347,460,1514,2327,3340,3940,6154,6220,7022,9100,9338,10152,11972,11980,13090,14500,14860,
12,148,348,461,1515,2328,3341,3941,6155,6221,7023,9101,9339,10153,11973,11981,13091,14501,14861,
13,149,349,462,1516,2329,3342,3942,6156,6222,7024,9102,9340,10154,11974,11982,13092,14502,14862,
14,150,350,463,1517,2330,3343,3943,6157,6223,7025,9103,9341,10155,11975,11983,13093,14503,14863,
15,151,351,464,1518,2331,3344,3944,6158,6224,7026,9104,9342,10156,11976,11984,13094,14504,14864,
16,152,352,465,1519,2332,3345,3945,6159,6225,7027,9105,9343,10157,11977,11985,13095,14505,14865,
17,153,353,466,1520,2333,3346,3946,6160,6226,7028,9106,9344,10158,11978,11986,13096,14506,14866,
18,154,354,467,1521,2334,3347,3947,6161,6227,7029,9107,9345,10159,11979,11987,13097,14507,14867,
19,155,355,468,1522,2335,3348,3948,6162,6228,7030,9108,9346,10160,11980,11988,13098,14508,14868,
20,156,356,469,1523,2336,3349,3949,6163,6229,7031,9109,9347,10161,11981,11989,13099,14509,14869,
21,157,357,470,1524,2337,3350,3950,6164,6230,7032,9110,9348,10162,11982,11990,13100,14510,14870,
22,158,358,471,1525,2338,3351,3951,6165,6231,7033,9111,9349,10163,11983,11991,13101,14511,14871,
23,159,359,472,1526,2339,3352,3952,6166,6232,7034,9112,9350,10164,11984,11992,13102,14512,14872,
0,24,160,473,1527,2340,3353,3953,6167,6233,7035,9113,9351,10165,11985,11993,13103,14513,14873,
1,25,161,474,1528,2341,3354,3954,6168,6234,7036,9114,9352,10166,11986,11994,13104,14514,14874,
2,26,162,475,1529,2342,3355,3955,6169,6235,7037,9115,9353,10167,11987,11995,13105,14515,14875,
3,27,163,476,1530,2343,3356,3956,6170,6236,7038,9116,9354,10168,11988,11996,13106,14516,14876,
4,28,164,477,1531,2344,3357,3957,6171,6237,7039,9117,9355,10169,11989,11997,13107,14517,14877,
5,29,165,478,1532,2345,3358,3958,6172,6238,7040,9118,9356,10170,11990,11998,13108,14518,14878,
6,30,166,479,1533,2346,3359,3959,6173,6239,7041,9119,9357,10171,11991,11999,13109,14519,14879,
7,31,167,480,1534,2347,3360,3600,6174,6240,7042,9120,9358,10172,11992,12000,13110,14520,14880,
8,32,168,481,1535,2348,3361,3601,6175,6241,7043,9121,9359,10173,11993,12001,13111,14521,14881,
9,33,169,482,1536,2349,3362,3602,6176,6242,7044,9000,9122,10174,11994,12002,13112,14522,14882,
10,34,170,483,1537,2350,3363,3603,6177,6243,7045,9001,9123,10175,11995,12003,13113,14523,14883,
11,35,171,484,1538,2351,3364,3604,6178,6244,7046,9002,9124,10176,11996,12004,13114,14524,14884,
12,36,172,485,1539,2352,3365,3605,6179,6245,7047,9003,9125,10177,11997,12005,13115,14525,14885,
13,37,173,486,1540,2353,3366,3606,6180,6246,7048,9004,9126,10178,11998,12006,13116,14526,14886,
14,38,174,487,1541,2354,3367,3607,6181,6247,7049,9005,9127,10179,11999,12007,13117,14527,14887,
15,39,175,488,1542,2355,3368,3608,6182,6248,7050,9006,9128,10180,12000,12008,13118,14528,14888,
16,40,176,489,1543,2356,3369,3609,6183,6249,7051,9007,9129,10181,12001,12009,13119,14529,14889,
17,41,177,490,1544,2357,3370,3610,6184,6250,7052,9008,9130,10182,12002,12010,13120,14530,14890,
18,42,178,491,1545,2358,3371,3611,6185,6251,7053,9009,9131,10183,12003,12011,13121,14531,14891,
19,43,179,492,1546,2359,3372,3612,6186,6252,7054,9010,9132,10184,12004,12012,13122,14532,14892,
20,44,180,493,1547,2360,3373,3613,6187,6253,7055,9011,9133,10185,12005,12013,13123,14533,14893,
21,45,181,494,1548,2361,3374,3614,6188,6254,7056,9012,9134,10186,12006,12014,13124,14534,14894,
22,46,182,495,1549,2362,3375,3615,6189,6255,7057,9013,9135,10187,12007,12015,13125,14535,14895,
23,47,183,496,1550,2363,3376,3616,6190,6256,7058,9014,9136,10188,12008,12016,13126,14536,14896,
24,48,184,497,1551,2364,3377,3617,6191,6257,7059,9015,9137,10189,12009,12017,13127,14537,14897,
25,49,185,498,1552,2365,3378,3618,6192,6258,7060,9016,9138,10190,12010,12018,13128,14538,14898,
26,50,186,499,1553,2366,3379,3619,6193,6259,7061,9017,9139,10191,12011,12019,13129,14539,14899,
27,51,187,500,1554,2367,3380,3620,6194,6260,7062,9018,9140,10192,12012,12020,13130,14540,14900,
28,52,188,501,1555,2368,3381,3621,6195,6261,7063,9019,9141,10193,12013,12021,13131,14541,14901,
29,53,189,502,1556,2369,3382,3622,6196,6262,7064,9020,9142,10194,12014,12022,13132,14542,14902,
30,54,190,503,1557,2370,3383,3623,6197,6263,7065,9021,9143,10195,12015,12023,13133,14543,14903,
31,55,191,504,1558,2371,3384,3624,6198,6264,7066,9022,9144,10196,12016,12024,13134,14544,14904,
32,56,192,505,1559,2372,3385,3625,6199,6265,7067,9023,9145,10197,12017,12025,13135,14545,14905,
33,57,193,506,1560,2373,3386,3626,6200,6266,7068,9024,9146,10198,12018,12026,13136,14546,14906,
34,58,194,507,1561,2374,3387,3627,6201,6267,7069,9025,9147,10199,12019,12027,13137,14547,14907,
35,59,195,508,1562,2375,3388,3628,6202,6268,7070,9026,9148,10200,12020,12028,13138,14548,14908,
36,60,196,509,1563,2376,3389,3629,6203,6269,7071,9027,9149,10201,12021,12029,13139,14549,14909,
37,61,197,510,1564,2377,3390,3630,6204,6270,7072,9028,9150,10202,12022,12030,13140,14550,14910,
38,62,198,511,1565,2378,3391,3631,6205,6271,7073,9029,9151,10203,12023,12031,13141,14551,14911,
39,63,199,512,1566,2379,3392,3632,6206,6272,7074,9030,9152,10204,12024,12032,13142,14552,14912,
40,64,200,513,1567,2380,3393,3633,6207,6273,7075,9031,9153,10205,12025,12033,13143,14553,14913,
41,65,201,514,1568,2381,3394,3634,6208,6274,7076,9032,9154,10206,12026,12034,13144,14554,14914,
42,66,202,515,1569,2382,3395,3635,6209,6275,7077,9033,9155,10207,12027,12035,13145,14555,14915,
43,67,203,516,1570,2383,3396,3636,6210,6276,7078,9034,9156,10208,12028,12036,13146,14556,14916,
44,68,204,517,1571,2384,3397,3637,6211,6277,7079,9035,9157,10209,12029,12037,13147,14557,14917,
45,69,205,518,1572,2385,3398,3638,6212,6278,7080,9036,9158,10210,12030,12038,13148,14558,14918,
46,70,206,519,1573,2386,3399,3639,6213,6279,7081,9037,9159,10211,12031,12039,13149,14559,14919,
47,71,207,520,1574,2387,3400,3640,6214,6280,7082,9038,9160,10212,12032,12040,13150,14560,14920,
48,72,208,521,1575,2388,3401,3641,6215,6281,7083,9039,9161,10213,12033,12041,13151,14561,14921,
49,73,209,522,1576,2389,3402,3642,6216,6282,7084,9040,9162,10214,12034,12042,13152,14562,14922,
50,74,210,523,1577,2390,3403,3643,6217,6283,7085,9041,9163,10215,12035,12043,13153,14563,14923,
51,75,211,524,1578,2391,3404,3644,6218,6284,7086,9042,9164,10216,12036,12044,13154,14564,14924,
52,76,212,525,1579,2392,3405,3645,6219,6285,7087,9043,9165,10217,12037,12045,13155,14565,14925,
53,77,213,526,1580,2393,3406,3646,6220,6286,7088,9044,9166,10218,12038,12046,13156,14566,14926,
54,78,214,527,1581,2394,3407,3647,6221,6287,7089,9045,9167,10219,12039,12047,13157,14567,14927,
55,79,215,528,1582,2395,3408,3648,6222,6288,7090,9046,9168,10220,12040,12048,13158,14568,14928,
56,80,216,529,1583,2396,3409,3649,6223,6289,7091,9047,9169,10221,12041,12049,13159,14569,14929,
57,81,217,530,1584,2397,3410,3650,6224,6290,7092,9048,9170,10222,12042,12050,13160,14570,14930,
58,82,218,531,1585,2398,3411,3651,6225,6291,7093,9049,9171,10223,12043,12051,13161,14571,14931,
59,83,219,532,1586,2399,3412,3652,6226,6292,7094,9050,9172,10224,12044,12052,13162,14572,14932,
60,84,220,533,1587,2400,3413,3653,6227,6293,7095,9051,9173,10225,12045,12053,13163,14573,14933,
61,85,221,534,1588,2401,3414,3654,6228,6294,7096,9052,9174,10226,12046,12054,13164,14574,14934,
62,86,222,535,1589,2402,3415,3655,6229,6295,7097,9053,9175,10227,12047,12055,13165,14575,14935,
63,87,223,536,1590,2403,3416,3656,6230,6296,7098,9054,9176,10228,12048,12056,13166,14576,14936,
64,88,224,537,1591,2404,3417,3657,6231,6297,7099,9055,9177,10229,12049,12057,13167,14577,14937,
65,89,225,538,1592,2405,3418,3658,6232,6298,7100,9056,9178,10230,12050,12058,13168,14578,14938,
66,90,226,539,1593,2406,3419,3659,6233,6299,7101,9057,9179,10231,12051,12059,13169,14579,14939,
67,91,227,540,1594,2407,3420,3660,6234,6300,7102,9058,9180,10232,12052,12060,13170,14580,14940,
68,92,228,541,1595,2408,3421,3661,6235,6301,7103,9059,9181,10233,12053,12061,13171,14581,14941,
69,93,229,542,1596,2409,3422,3662,6236,6302,7104,9060,9182,10234,12054,12062,13172,14582,14942,
70,94,230,543,1597,2410,3423,3663,6237,6303,7105,9061,9183,10235,12055,12063,13173,14583,14943,
71,95,231,544,1598,2411,3424,3664,6238,6304,7106,9062,9184,10236,12056,12064,13174,14584,14944,
72,96,232,545,1599,2412,3425,3665,6239,6305,7107,9063,9185,10237,12057,12065,13175,14585,14945,
73,97,233,546,1600,2413,3426,3666,6240,6306,7108,9064,9186,10238,12058,12066,13176,14586,14946,
74,98,234,547,1601,2414,3427,3667,6241,6307,7109,9065,9187,10239,12059,12067,13177,14587,14947,
75,99,235,548,1602,2415,3428,3668,6242,6308,7110,9066,9188,10240,12060,12068,13178,14588,14948,
76,100,236,549,1603,2416,3429,3669,6243,6309,7111,9067,9189,10241,12061,12069,13179,14589,14949,
77,101,237,550,1604,2417,3430,3670,6244,6310,7112,9068,9190,10242,12062,12070,13180,14590,14950,
78,102,238,551,1605,2418,3431,3671,6245,6311,7113,9069,9191,10243,12063,12071,13181,14591,14951,
79,103,239,552,1606,2419,3432,3672,6246,6312,7114,9070,9192,10244,12064,12072,13182,14592,14952,
80,104,240,553,1607,2420,3433,3673,6247,6313,7115,9071,9193,10245,12065,12073,13183,14593,14953,
81,105,241,554,1608,2421,3434,3674,6248,6314,7116,9072,9194,10246,12066,12074,13184,14594,14954,
82,106,242,555,1609,2422,3435,3675,6249,6315,7117,9073,9195,10247,12067,12075,13185,14595,14955,
83,107,243,556,1610,2423,3436,3676,6250,6316,7118,9074,9196,10248,12068,12076,13186,14596,14956,
84,108,244,557,1611,2424,3437,3677,6251,6317,7119,9075,9197,10249,12069,12077,13187,14597,14957,
85,109,245,558,1612,2425,3438,3678,6252,6318,7120,9076,9198,10250,12070,12078,13188,14598,14958,
86,110,246,559,1613,2426,3439,3679,6253,6319,7121,9077,9199,10251,12071,12079,13189,14599,14959,
87,111,247,560,1614,2427,3440,3680,6254,6320,7122,9078,9200,10252,12072,12080,13190,14600,14960,
88,112,248,561,1615,2428,3441,3681,6255,6321,7123,9079,9201,10253,12073,12081,13191,14601,14961,
89,113,249,562,1616,2429,3442,3682,6256,6322,7124,9080,9202,10254,12074,12082,13192,14602,14962,
90,114,250,563,1617,2430,3443,3683,6257,6323,7125,9081,9203,10255,12075,12083,13193,14603,14963,
91,115,251,564,1618,2431,3444,3684,6258,6324,7126,9082,9204,10256,12076,12084,13194,14604,14964,
92,116,252,565,1619,2432,3445,3685,6259,6325,7127,9083,9205,10257,12077,12085,13195,14605,14965,
93,117,253,566,1620,2433,3446,3686,6260,6326,7128,9084,9206,10258,12078,12086,13196,14606,14966,
94,118,254,567,1621,2434,3447,3687,6261,6327,7129,9085,9207,10259,12079,12087,13197,14607,14967,
95,119,255,568,1622,2435,3448,3688,6262,6328,7130,9086,9208,10260,12080,12088,13198,14608,14968,
96,120,256,569,1623,2436,3449,3689,6263,6329,7131,9087,9209,10261,12081,12089,13199,14609,14969,
97,121,257,570,1624,2437,3450,3690,6264,6330,7132,9088,9210,10262,12082,12090,13200,14610,14970,
98,122,258,571,1625,2438,3451,3691,6265,6331,7133,9089,9211,10263,12083,12091,13201,14611,14971,
99,123,259,572,1626,2439,3452,3692,6266,6332,7134,9090,9212,10264,12084,12092,13202,14612,14972,
100,124,260,573,1627,2440,3453,3693,6267,6333,7135,9091,9213,10265,12085,12093,13203,14613,14973,
101,125,261,574,1628,2441,3454,3694,6268,6334,7136,9092,9214,10266,12086,12094,13204,14614,14974,
102,126,262,575,1629,2442,3455,3695,6269,6335,7137,9093,9215,10267,12087,12095,13205,14615,14975,
103,127,263,576,1630,2443,3456,3696,6270,6336,7138,9094,9216,10268,12088,12096,13206,14616,14976,
104,128,264,577,1631,2444,3457,3697,6271,6337,7139,9095,9217,10269,12089,12097,13207,14617,14977,
105,129,265,578,1632,2445,3458,3698,6272,6338,7140,9096,9218,10270,12090,12098,13208,14618,14978,
106,130,266,579,1633,2446,3459,3699,6273,6339,7141,9097,9219,10271,12091,12099,13209,14619,14979,
107,131,267,580,1634,2447,3460,3700,6274,6340,7142,9098,9220,10272,12092,12100,13210,14620,14980,
108,132,268,581,1635,2448,3461,3701,6275,6341,7143,9099,9221,10273,12093,12101,13211,14621,14981,
109,133,269,582,1636,2449,3462,3702,6276,6342,7144,9100,9222,10274,12094,12102,13212,14622,14982,
110,134,270,583,1637,2450,3463,3703,6277,6343,7145,9101,9223,10275,12095,12103,13213,14623,14983,
111,135,271,584,1638,2451,3464,3704,6278,6344,7146,9102,9224,10276,12096,12104,13214,14624,14984,
112,136,272,585,1639,2452,3465,3705,6279,6345,7147,9103,9225,10277,12097,12105,13215,14625,14985,
113,137,273,586,1640,2453,3466,3706,6280,6346,7148,9104,9226,10278,12098,12106,13216,14626,14986,
114,138,274,587,1641,2454,3467,3707,6281,6347,7149,9105,9227,10279,12099,12107,13217,14627,14987,
115,139,275,588,1642,2455,3468,3708,6282,6348,7150,9106,9228,10280,12100,12108,13218,14628,14988,
116,140,276,589,1643,2456,3469,3709,6283,6349,7151,9107,9229,10281,12101,12109,13219,14629,14989,
117,141,277,590,1644,2457,3470,3710,6284,6350,7152,9108,9230,10282,12102,12110,13220,14630,14990,
118,142,278,591,1645,2458,3471,3711,6285,6351,7153,9109,9231,10283,12103,12111,13221,14631,14991,
119,143,279,592,1646,2459,3472,3712,6286,6352,7154,9110,9232,10284,12104,12112,13222,14632,14992,
120,144,280,593,1647,2460,3473,3713,6287,6353,7155,9111,9233,10285,12105,12113,13223,14633,14993,
121,145,281,594,1648,2461,3474,3714,6288,6354,7156,9112,9234,10286,12106,12114,13224,14634,14994,
122,146,282,595,1649,2462,3475,3715,6289,6355,7157,9113,9235,10287,12107,12115,13225,14635,14995,
123,147,283,596,1650,2463,3476,3716,6290,6356,7158,9114,9236,10288,12108,12116,13226,14636,14996,
124,148,284,597,1651,2464,3477,3717,6291,6357,7159,9115,9237,10289,12109,12117,13227,14637,14997,
125,149,285,598,1652,2465,3478,3718,6292,6358,7160,9116,9238,10290,12110,12118,13228,14638,14998,
126,150,286,599,1653,2466,3479,3719,6293,6359,7161,9117,9239,10291,12111,12119,13229,14639,14999,
127,151,287,600,1654,2467,3480,3720,6294,6360,7162,9118,9240,10292,12112,12120,13230,14640,15000,
128,152,288,601,1655,2468,3481,3721,6295,6361,7163,9119,9241,10293,12113,12121,13231,14641,15001,
129,153,289,602,1656,2469,3482,3722,6296,6362,7164,9120,9242,10294,12114,12122,13232,14642,15002,
130,154,290,603,1657,2470,3483,3723,6297,6363,7165,9121,9243,10295,12115,12123,13233,14643,15003,
131,155,291,604,1658,2471,3484,3724,6298,6364,7166,9122,9244,10296,12116,12124,13234,14644,15004,
132,156,292,605,1659,2472,3485,3725,6299,6365,7167,9123,9245,10297,12117,12125,13235,14645,15005,
133,157,293,606,1660,2473,3486,3726,6300,6366,7168,9124,9246,10298,12118,12126,13236,14646,15006,
134,158,294,607,1661,2474,3487,3727,6301,6367,7169,9125,9247,10299,12119,12127,13237,14647,15007,
135,159,295,608,1662,2475,3488,3728,6302,6368,7170,9126,9248,10300,12120,12128,13238,14648,15008,
136,160,296,609,1663,2476,3489,3729,6303,6369,7171,9127,9249,10301,12121,12129,13239,14649,15009,
137,161,297,610,1664,2477,3490,3730,6304,6370,7172,9128,9250,10302,12122,12130,13240,14650,15010,
138,162,298,611,1665,2478,3491,3731,6305,6371,7173,9129,9251,10303,12123,12131,13241,14651,15011,
139,163,299,612,1666,2479,3492,3732,6306,6372,7174,9130,9252,10304,12124,12132,13242,14652,15012,
140,164,300,613,1667,2480,3493,3733,6307,6373,7175,9131,9253,10305,12125,12133,13243,14653,15013,
141,165,301,614,1668,2481,3494,3734,6308,6374,7176,9132,9254,10306,12126,12134,13244,14654,15014,
142,166,302,615,1669,2482,3495,3735,6309,6375,7177,9133,9255,10307,12127,12135,13245,14655,15015,
143,167,303,616,1670,2483,3496,3736,6310,6376,7178,9134,9256,10308,12128,12136,13246,14656,15016,
144,168,304,617,1671,2484,3497,3737,6311,6377,7179,9135,9257,10309,12129,12137,13247,14657,15017,
145,169,305,618,1672,2485,3498,3738,6312,6378,7180,9136,9258,10310,12130,12138,13248,14658,15018,
146,170,306,619,1673,2486,3499,3739,6313,6379,7181,9137,9259,10311,12131,12139,13249,14659,15019,
147,171,307,620,1674,2487,3500,3740,6314,6380,7182,9138,9260,10312,12132,12140,13250,14660,15020,
148,172,308,621,1675,2488,3501,3741,6315,6381,7183,9139,9261,10313,12133,12141,13251,14661,15021,
149,173,309,622,1676,2489,3502,3742,6316,6382,7184,9140,9262,10314,12134,12142,13252,14662,15022,
150,174,310,623,1677,2490,3503,3743,6317,6383,7185,9141,9263,10315,12135,12143,13253,14663,15023,
151,175,311,624,1678,2491,3504,3744,6318,6384,7186,9142,9264,10316,12136,12144,13254,14664,15024,
152,176,312,625,1679,2492,3505,3745,6319,6385,7187,9143,9265,10317,12137,12145,13255,14665,15025,
153,177,313,626,1680,2493,3506,3746,6320,6386,7188,9144,9266,10318,12138,12146,13256,14666,15026,
154,178,314,627,1681,2494,3507,3747,6321,6387,7189,9145,9267,10319,12139,12147,13257,14667,15027,
155,179,315,628,1682,2495,3508,3748,6322,6388,7190,9146,9268,10320,12140,12148,13258,14668,15028,
156,180,316,629,1683,2496,3509,3749,6323,6389,7191,9147,9269,10321,12141,12149,13259,14669,15029,
157,181,317,630,1684,2497,3510,3750,6324,6390,7192,9148,9270,10322,12142,12150,13260,14670,15030,
158,182,318,631,1685,2498,3511,3751,6325,6391,7193,9149,9271,10323,12143,12151,13261,14671,15031,
159,183,319,632,1686,2499,3512,3752,6326,6392,7194,9150,9272,10324,12144,12152,13262,14672,15032,
160,184,320,633,1687,2500,3513,3753,6327,6393,7195,9151,9273,10325,12145,12153,13263,14673,15033,
161,185,321,634,1688,2501,3514,3754,6328,6394,7196,9152,9274,10326,12146,12154,13264,14674,15034,
162,186,322,635,1689,2502,3515,3755,6329,6395,7197,9153,9275,10327,12147,12155,13265,14675,15035,
163,187,323,636,1690,2503,3516,3756,6330,6396,7198,9154,9276,10328,12148,12156,13266,14676,15036,
164,188,324,637,1691,2504,3517,3757,6331,6397,7199,9155,9277,10329,12149,12157,13267,14677,15037,
165,189,325,638,1692,2505,3518,3758,6332,6398,6840,9156,9278,10330,12150,12158,13268,14678,15038,
166,190,326,639,1693,2506,3519,3759,6333,6399,6841,9157,9279,10331,12151,12159,13269,14679,15039,
167,191,327,640,1694,2507,3520,3760,6334,6400,6842,9158,9280,10332,12152,12160,13270,14680,15040,
168,192,328,641,1695,2508,3521,3761,6335,6401,6843,9159,9281,10333,12153,12161,13271,14681,15041,
169,193,329,642,1696,2509,3522,3762,6336,6402,6844,9160,9282,10334,12154,12162,13272,14682,15042,
170,194,330,643,1697,2510,3523,3763,6337,6403,6845,9161,9283,10335,12155,12163,13273,14683,15043,
171,195,331,644,1698,2511,3524,3764,6338,6404,6846,9162,9284,10336,12156,12164,13274,14684,15044,
172,196,332,645,1699,2512,3525,3765,6339,6405,6847,9163,9285,10337,12157,12165,13275,14685,15045,
173,197,333,646,1700,2513,3526,3766,6340,6406,6848,9164,9286,10338,12158,12166,13276,14686,15046,
174,198,334,647,1701,2514,3527,3767,6341,6407,6849,9165,9287,10339,12159,12167,13277,14687,15047,
175,199,335,648,1702,2515,3528,3768,6342,6408,6850,9166,9288,10340,12160,12168,13278,14688,15048,
176,200,336,649,1703,2516,3529,3769,6343,6409,6851,9167,9289,10341,12161,12169,13279,14689,15049,
177,201,337,650,1704,2517,3530,3770,6344,6410,6852,9168,9290,10342,12162,12170,13280,14690,15050,
178,202,338,651,1705,2518,3531,3771,6345,6411,6853,9169,9291,10343,12163,12171,13281,14691,15051,
179,203,339,652,1706,2519,3532,3772,6346,6412,6854,9170,9292,10344,12164,12172,13282,14692,15052,
180,204,340,653,1707,2160,3533,3773,6347,6413,6855,9171,9293,10345,12165,12173,13283,14693,15053,
181,205,341,654,1708,2161,3534,3774,6348,6414,6856,9172,9294,10346,12166,12174,13284,14694,15054,
182,206,342,655,1709,2162,3535,3775,6349,6415,6857,9173,9295,10347,12167,12175,13285,14695,15055,
183,207,343,656,1710,2163,3536,3776,6350,6416,6858,9174,9296,10348,12168,12176,13286,14696,15056,
184,208,344,657,1711,2164,3537,3777,6351,6417,6859,9175,9297,10349,12169,12177,13287,14697,15057,
185,209,345,658,1712,2165,3538,3778,6352,6418,6860,9176,9298,10350,12170,12178,13288,14698,15058,
186,210,346,659,1713,2166,3539,3779,6353,6419,6861,9177,9299,10351,12171,12179,13289,14699,15059,
187,211,347,660,1714,2167,3540,3780,6354,6420,6862,9178,9300,10352,12172,12180,13290,14700,15060,
188,212,348,661,1715,2168,3541,3781,6355,6421,6863,9179,9301,10353,12173,12181,13291,14701,15061,
189,213,349,662,1716,2169,3542,3782,6356,6422,6864,9180,9302,10354,12174,12182,13292,14702,15062,
190,214,350,663,1717,2170,3543,3783,6357,6423,6865,9181,9303,10355,12175,12183,13293,14703,15063,
191,215,351,664,1718,2171,3544,3784,6358,6424,6866,9182,9304,10356,12176,12184,13294,14704,15064,
192,216,352,665,1719,2172,3545,3785,6359,6425,6867,9183,9305,10357,12177,12185,13295,14705,15065,
193,217,353,666,1720,2173,3546,3786,6360,6426,6868,9184,9306,10358,12178,12186,13296,14706,15066,
194,218,354,667,1721,2174,3547,3787,6361,6427,6869,9185,9307,10359,12179,12187,13297,14707,15067,
195,219,355,668,1722,2175,3548,3788,6362,6428,6870,9186,9308,10360,12180,12188,13298,14708,15068,
196,220,356,669,1723,2176,3549,3789,6363,6429,6871,9187,9309,10361,12181,12189,13299,14709,15069,
197,221,357,670,1724,2177,3550,3790,6364,6430,6872,9188,9310,10362,12182,12190,13300,14710,15070,
198,222,358,671,1725,2178,3551,3791,6365,6431,6873,9189,9311,10363,12183,12191,13301,14711,15071,
199,223,359,672,1726,2179,3552,3792,6366,6432,6874,9190,9312,10364,12184,12192,13302,14712,15072,
0,200,224,673,1727,2180,3553,3793,6367,6433,6875,9191,9313,10365,12185,12193,13303,14713,15073,
1,201,225,674,1728,2181,3554,3794,6368,6434,6876,9192,9314,10366,12186,12194,13304,14714,15074,
2,202,226,675,1729,2182,3555,3795,6369,6435,6877,9193,9315,10367,12187,12195,13305,14715,15075,
3,203,227,676,1730,2183,3556,3796,6370,6436,6878,9194,9316,10368,12188,12196,13306,14716,15076,
4,204,228,677,1731,2184,3557,3797,6371,6437,6879,9195,9317,10369,12189,12197,13307,14717,15077,
5,205,229,678,1732,2185,3558,3798,6372,6438,6880,9196,9318,10370,12190,12198,13308,14718,15078,
6,206,230,679,1733,2186,3559,3799,6373,6439,6881,9197,9319,10371,12191,12199,13309,14719,15079,
7,207,231,680,1734,2187,3560,3800,6374,6440,6882,9198,9320,10372,12192,12200,13310,14720,15080,
8,208,232,681,1735,2188,3561,3801,6375,6441,6883,9199,9321,10373,12193,12201,13311,14721,15081,
9,209,233,682,1736,2189,3562,3802,6376,6442,6884,9200,9322,10374,12194,12202,13312,14722,15082,
10,210,234,683,1737,2190,3563,3803,6377,6443,6885,9201,9323,10375,12195,12203,13313,14723,15083,
11,211,235,684,1738,2191,3564,3804,6378,6444,6886,9202,9324,10376,12196,12204,13314,14724,15084,
12,212,236,685,1739,2192,3565,3805,6379,6445,6887,9203,9325,10377,12197,12205,13315,14725,15085,
13,213,237,686,1740,2193,3566,3806,6380,6446,6888,9204,9326,10378,12198,12206,13316,14726,15086,
14,214,238,687,1741,2194,3567,3807,6381,6447,6889,9205,9327,10379,12199,12207,13317,14727,15087,
15,215,239,688,1742,2195,3568,3808,6382,6448,6890,9206,9328,10380,12200,12208,13318,14728,15088,
16,216,240,689,1743,2196,3569,3809,6383,6449,6891,9207,9329,10381,12201,12209,13319,14729,15089,
17,217,241,690,1744,2197,3570,3810,6384,6450,6892,9208,9330,10382,12202,12210,12960,14730,15090,
18,218,242,691,1745,2198,3571,3811,6385,6451,6893,9209,9331,10383,12203,12211,12961,14731,15091,
19,219,243,692,1746,2199,3572,3812,6386,6452,6894,9210,9332,10384,12204,12212,12962,14732,15092,
20,220,244,693,1747,2200,3573,3813,6387,6453,6895,9211,9333,10385,12205,12213,12963,14733,15093,
21,221,245,694,1748,2201,3574,3814,6388,6454,6896,9212,9334,10386,12206,12214,12964,14734,15094,
22,222,246,695,1749,2202,3575,3815,6389,6455,6897,9213,9335,10387,12207,12215,12965,14735,15095,
23,223,247,696,1750,2203,3576,3816,6390,6456,6898,9214,9336,10388,12208,12216,12966,14736,15096,
24,224,248,697,1751,2204,3577,3817,6391,6457,6899,9215,9337,10389,12209,12217,12967,14737,15097,
25,225,249,698,1752,2205,3578,3818,6392,6458,6900,9216,9338,10390,12210,12218,12968,14738,15098,
26,226,250,699,1753,2206,3579,3819,6393,6459,6901,9217,9339,10391,12211,12219,12969,14739,15099,
27,227,251,700,1754,2207,3580,3820,6394,6460,6902,9218,9340,10392,12212,12220,12970,14740,15100,
28,228,252,701,1755,2208,3581,3821,6395,6461,6903,9219,9341,10393,12213,12221,12971,14741,15101,
29,229,253,702,1756,2209,3582,3822,6396,6462,6904,9220,9342,10394,12214,12222,12972,14742,15102,
30,230,254,703,1757,2210,3583,3823,6397,6463,6905,9221,9343,10395,12215,12223,12973,14743,15103,
31,231,255,704,1758,2211,3584,3824,6398,6464,6906,9222,9344,10396,12216,12224,12974,14744,15104,
32,232,256,705,1759,2212,3585,3825,6399,6465,6907,9223,9345,10397,12217,12225,12975,14745,15105,
33,233,257,706,1760,2213,3586,3826,6400,6466,6908,9224,9346,10398,12218,12226,12976,14746,15106,
34,234,258,707,1761,2214,3587,3827,6401,6467,6909,9225,9347,10399,12219,12227,12977,14747,15107,
35,235,259,708,1762,2215,3588,3828,6402,6468,6910,9226,9348,10400,12220,12228,12978,14748,15108,
36,236,260,709,1763,2216,3589,3829,6403,6469,6911,9227,9349,10401,12221,12229,12979,14749,15109,
37,237,261,710,1764,2217,3590,3830,6404,6470,6912,9228,9350,10402,12222,12230,12980,14750,15110,
38,238,262,711,1765,2218,3591,3831,6405,6471,6913,9229,9351,10403,12223,12231,12981,14751,15111,
39,239,263,712,1766,2219,3592,3832,6406,6472,6914,9230,9352,10404,12224,12232,12982,14752,15112,
40,240,264,713,1767,2220,3593,3833,6407,6473,6915,9231,9353,10405,12225,12233,12983,14753,15113,
41,241,265,714,1768,2221,3594,3834,6408,6474,6916,9232,9354,10406,12226,12234,12984,14754,15114,
42,242,266,715,1769,2222,3595,3835,6409,6475,6917,9233,9355,10407,12227,12235,12985,14755,15115,
43,243,267,716,1770,2223,3596,3836,6410,6476,6918,9234,9356,10408,12228,12236,12986,14756,15116,
44,244,268,717,1771,2224,3597,3837,6411,6477,6919,9235,9357,10409,12229,12237,12987,14757,15117,
45,245,269,718,1772,2225,3598,3838,6412,6478,6920,9236,9358,10410,12230,12238,12988,14758,15118,
46,246,270,719,1773,2226,3599,3839,6413,6479,6921,9237,9359,10411,12231,12239,12989,14759,15119,
10,319,720,1729,3388,3600,4019,4843,4885,6480,8123,8141,9360,10565,12240,12880,14760,15120,
11,320,721,1730,3389,3601,4020,4844,4886,6481,8124,8142,9361,10566,12241,12881,14761,15121,
12,321,722,1731,3390,3602,4021,4845,4887,6482,8125,8143,9362,10567,12242,12882,14762,15122,
13,322,723,1732,3391,3603,4022,4846,4888,6483,8126,8144,9363,10568,12243,12883,14763,15123,
14,323,724,1733,3392,3604,4023,4847,4889,6484,8127,8145,9364,10569,12244,12884,14764,15124,
15,324,725,1734,3393,3605,4024,4848,4890,6485,8128,8146,9365,10570,12245,12885,14765,15125,
16,325,726,1735,3394,3606,4025,4849,4891,6486,8129,8147,9366,10571,12246,12886,14766,15126,
17,326,727,1736,3395,3607,4026,4850,4892,6487,8130,8148,9367,10572,12247,12887,14767,15127,
18,327,728,1737,3396,3608,4027,4851,4893,6488,8131,8149,9368,10573,12248,12888,14768,15128,
19,328,729,1738,3397,3609,4028,4852,4894,6489,8132,8150,9369,10574,12249,12889,14769,15129,
20,329,730,1739,3398,3610,4029,4853,4895,6490,8133,8151,9370,10575,12250,12890,14770,15130,
21,330,731,1740,3399,3611,4030,4854,4896,6491,8134,8152,9371,10576,12251,12891,14771,15131,
22,331,732,1741,3400,3612,4031,4855,4897,6492,8135,8153,9372,10577,12252,12892,14772,15132,
23,332,733,1742,3401,3613,4032,4856,4898,6493,8136,8154,9373,10578,12253,12893,14773,15133,
24,333,734,1743,3402,3614,4033,4857,4899,6494,8137,8155,9374,10579,12254,12894,14774,15134,
25,334,735,1744,3403,3615,4034,4858,4900,6495,8138,8156,9375,10580,12255,12895,14775,15135,
26,335,736,1745,3404,3616,4035,4859,4901,6496,8139,8157,9376,10581,12256,12896,14776,15136,
27,336,737,1746,3405,3617,4036,4860,4902,6497,8140,8158,9377,10582,12257,12897,14777,15137,
28,337,738,1747,3406,3618,4037,4861,4903,6498,8141,8159,9378,10583,12258,12898,14778,15138,
29,338,739,1748,3407,3619,4038,4862,4904,6499,8142,8160,9379,10584,12259,12899,14779,15139,
30,339,740,1749,3408,3620,4039,4863,4905,6500,8143,8161,9380,10585,12260,12900,14780,15140,
31,340,741,1750,3409,3621,4040,4864,4906,6501,8144,8162,9381,10586,12261,12901,14781,15141,
32,341,742,1751,3410,3622,4041,4865,4907,6502,8145,8163,9382,10587,12262,12902,14782,15142,
33,342,743,1752,3411,3623,4042,4866,4908,6503,8146,8164,9383,10588,12263,12903,14783,15143,
34,343,744,1753,3412,3624,4043,4867,4909,6504,8147,8165,9384,10589,12264,12904,14784,15144,
35,344,745,1754,3413,3625,4044,4868,4910,6505,8148,8166,9385,10590,12265,12905,14785,15145,
36,345,746,1755,3414,3626,4045,4869,4911,6506,8149,8167,9386,10591,12266,12906,14786,15146,
37,346,747,1756,3415,3627,4046,4870,4912,6507,8150,8168,9387,10592,12267,12907,14787,15147,
38,347,748,1757,3416,3628,4047,4871,4913,6508,8151,8169,9388,10593,12268,12908,14788,15148,
39,348,749,1758,3417,3629,4048,4872,4914,6509,8152,8170,9389,10594,12269,12909,14789,15149,
40,349,750,1759,3418,3630,4049,4873,4915,6510,8153,8171,9390,10595,12270,12910,14790,15150,
41,350,751,1760,3419,3631,4050,4874,4916,6511,8154,8172,9391,10596,12271,12911,14791,15151,
42,351,752,1761,3420,3632,4051,4875,4917,6512,8155,8173,9392,10597,12272,12912,14792,15152,
43,352,753,1762,3421,3633,4052,4876,4918,6513,8156,8174,9393,10598,12273,12913,14793,15153,
44,353,754,1763,3422,3634,4053,4877,4919,6514,8157,8175,9394,10599,12274,12914,14794,15154,
45,354,755,1764,3423,3635,4054,4878,4920,6515,8158,8176,9395,10600,12275,12915,14795,15155,
46,355,756,1765,3424,3636,4055,4879,4921,6516,8159,8177,9396,10601,12276,12916,14796,15156,
47,356,757,1766,3425,3637,4056,4880,4922,6517,8160,8178,9397,10602,12277,12917,14797,15157,
48,357,758,1767,3426,3638,4057,4881,4923,6518,8161,8179,9398,10603,12278,12918,14798,15158,
49,358,759,1768,3427,3639,4058,4882,4924,6519,8162,8180,9399,10604,12279,12919,14799,15159,
50,359,760,1769,3428,3640,4059,4883,4925,6520,8163,8181,9400,10605,12280,12920,14800,15160,
0,51,761,1770,3429,3641,4060,4884,4926,6521,8164,8182,9401,10606,12281,12921,14801,15161,
1,52,762,1771,3430,3642,4061,4885,4927,6522,8165,8183,9402,10607,12282,12922,14802,15162,
2,53,763,1772,3431,3643,4062,4886,4928,6523,8166,8184,9403,10608,12283,12923,14803,15163,
3,54,764,1773,3432,3644,4063,4887,4929,6524,8167,8185,9404,10609,12284,12924,14804,15164,
4,55,765,1774,3433,3645,4064,4888,4930,6525,8168,8186,9405,10610,12285,12925,14805,15165,
5,56,766,1775,3434,3646,4065,4889,4931,6526,8169,8187,9406,10611,12286,12926,14806,15166,
6,57,767,1776,3435,3647,4066,4890,4932,6527,8170,8188,9407,10612,12287,12927,14807,15167,
7,58,768,1777,3436,3648,4067,4891,4933,6528,8171,8189,9408,10613,12288,12928,14808,15168,
8,59,769,1778,3437,3649,4068,4892,4934,6529,8172,8190,9409,10614,12289,12929,14809,15169,
9,60,770,1779,3438,3650,4069,4893,4935,6530,8173,8191,9410,10615,12290,12930,14810,15170,
10,61,771,1780,3439,3651,4070,4894,4936,6531,8174,8192,9411,10616,12291,12931,14811,15171,
11,62,772,1781,3440,3652,4071,4895,4937,6532,8175,8193,9412,10617,12292,12932,14812,15172,
12,63,773,1782,3441,3653,4072,4896,4938,6533,8176,8194,9413,10618,12293,12933,14813,15173,
13,64,774,1783,3442,3654,4073,4897,4939,6534,8177,8195,9414,10619,12294,12934,14814,15174,
14,65,775,1784,3443,3655,4074,4898,4940,6535,8178,8196,9415,10620,12295,12935,14815,15175,
15,66,776,1785,3444,3656,4075,4899,4941,6536,8179,8197,9416,10621,12296,12936,14816,15176,
16,67,777,1786,3445,3657,4076,4900,4942,6537,8180,8198,9417,10622,12297,12937,14817,15177,
17,68,778,1787,3446,3658,4077,4901,4943,6538,8181,8199,9418,10623,12298,12938,14818,15178,
18,69,779,1788,3447,3659,4078,4902,4944,6539,8182,8200,9419,10624,12299,12939,14819,15179,
19,70,780,1789,3448,3660,4079,4903,4945,6540,8183,8201,9420,10625,12300,12940,14820,15180,
20,71,781,1790,3449,3661,4080,4904,4946,6541,8184,8202,9421,10626,12301,12941,14821,15181,
21,72,782,1791,3450,3662,4081,4905,4947,6542,8185,8203,9422,10627,12302,12942,14822,15182,
22,73,783,1792,3451,3663,4082,4906,4948,6543,8186,8204,9423,10628,12303,12943,14823,15183,
23,74,784,1793,3452,3664,4083,4907,4949,6544,8187,8205,9424,10629,12304,12944,14824,15184,
24,75,785,1794,3453,3665,4084,4908,4950,6545,8188,8206,9425,10630,12305,12945,14825,15185,
25,76,786,1795,3454,3666,4085,4909,4951,6546,8189,8207,9426,10631,12306,12946,14826,15186,
26,77,787,1796,3455,3667,4086,4910,4952,6547,8190,8208,9427,10632,12307,12947,14827,15187,
27,78,788,1797,3456,3668,4087,4911,4953,6548,8191,8209,9428,10633,12308,12948,14828,15188,
28,79,789,1798,3457,3669,4088,4912,4954,6549,8192,8210,9429,10634,12309,12949,14829,15189,
29,80,790,1799,3458,3670,4089,4913,4955,6550,8193,8211,9430,10635,12310,12950,14830,15190,
30,81,791,1440,3459,3671,4090,4914,4956,6551,8194,8212,9431,10636,12311,12951,14831,15191,
31,82,792,1441,3460,3672,4091,4915,4957,6552,8195,8213,9432,10637,12312,12952,14832,15192,
32,83,793,1442,3461,3673,4092,4916,4958,6553,8196,8214,9433,10638,12313,12953,14833,15193,
33,84,794,1443,3462,3674,4093,4917,4959,6554,8197,8215,9434,10639,12314,12954,14834,15194,
34,85,795,1444,3463,3675,4094,4918,4960,6555,8198,8216,9435,10640,12315,12955,14835,15195,
35,86,796,1445,3464,3676,4095,4919,4961,6556,8199,8217,9436,10641,12316,12956,14836,15196,
36,87,797,1446,3465,3677,4096,4920,4962,6557,8200,8218,9437,10642,12317,12957,14837,15197,
37,88,798,1447,3466,3678,4097,4921,4963,6558,8201,8219,9438,10643,12318,12958,14838,15198,
38,89,799,1448,3467,3679,4098,4922,4964,6559,8202,8220,9439,10644,12319,12959,14839,15199,
39,90,800,1449,3468,3680,4099,4923,4965,6560,8203,8221,9440,10645,12320,12600,14840,15200,
40,91,801,1450,3469,3681,4100,4924,4966,6561,8204,8222,9441,10646,12321,12601,14841,15201,
41,92,802,1451,3470,3682,4101,4925,4967,6562,8205,8223,9442,10647,12322,12602,14842,15202,
42,93,803,1452,3471,3683,4102,4926,4968,6563,8206,8224,9443,10648,12323,12603,14843,15203,
43,94,804,1453,3472,3684,4103,4927,4969,6564,8207,8225,9444,10649,12324,12604,14844,15204,
44,95,805,1454,3473,3685,4104,4928,4970,6565,8208,8226,9445,10650,12325,12605,14845,15205,
45,96,806,1455,3474,3686,4105,4929,4971,6566,8209,8227,9446,10651,12326,12606,14846,15206,
46,97,807,1456,3475,3687,4106,4930,4972,6567,8210,8228,9447,10652,12327,12607,14847,15207,
47,98,808,1457,3476,3688,4107,4931,4973,6568,8211,8229,9448,10653,12328,12608,14848,15208,
48,99,809,1458,3477,3689,4108,4932,4974,6569,8212,8230,9449,10654,12329,12609,14849,15209,
49,100,810,1459,3478,3690,4109,4933,4975,6570,8213,8231,9450,10655,12330,12610,14850,15210,
50,101,811,1460,3479,3691,4110,4934,4976,6571,8214,8232,9451,10656,12331,12611,14851,15211,
51,102,812,1461,3480,3692,4111,4935,4977,6572,8215,8233,9452,10657,12332,12612,14852,15212,
52,103,813,1462,3481,3693,4112,4936,4978,6573,8216,8234,9453,10658,12333,12613,14853,15213,
53,104,814,1463,3482,3694,4113,4937,4979,6574,8217,8235,9454,10659,12334,12614,14854,15214,
54,105,815,1464,3483,3695,4114,4938,4980,6575,8218,8236,9455,10660,12335,12615,14855,15215,
55,106,816,1465,3484,3696,4115,4939,4981,6576,8219,8237,9456,10661,12336,12616,14856,15216,
56,107,817,1466,3485,3697,4116,4940,4982,6577,8220,8238,9457,10662,12337,12617,14857,15217,
57,108,818,1467,3486,3698,4117,4941,4983,6578,8221,8239,9458,10663,12338,12618,14858,15218,
58,109,819,1468,3487,3699,4118,4942,4984,6579,8222,8240,9459,10664,12339,12619,14859,15219,
59,110,820,1469,3488,3700,4119,4943,4985,6580,8223,8241,9460,10665,12340,12620,14860,15220,
60,111,821,1470,3489,3701,4120,4944,4986,6581,8224,8242,9461,10666,12341,12621,14861,15221,
61,112,822,1471,3490,3702,4121,4945,4987,6582,8225,8243,9462,10667,12342,12622,14862,15222,
62,113,823,1472,3491,3703,4122,4946,4988,6583,8226,8244,9463,10668,12343,12623,14863,15223,
63,114,824,1473,3492,3704,4123,4947,4989,6584,8227,8245,9464,10669,12344,12624,14864,15224,
64,115,825,1474,3493,3705,4124,4948,4990,6585,8228,8246,9465,10670,12345,12625,14865,15225,
65,116,826,1475,3494,3706,4125,4949,4991,6586,8229,8247,9466,10671,12346,12626,14866,15226,
66,117,827,1476,3495,3707,4126,4950,4992,6587,8230,8248,9467,10672,12347,12627,14867,15227,
67,118,828,1477,3496,3708,4127,4951,4993,6588,8231,8249,9468,10673,12348,12628,14868,15228,
68,119,829,1478,3497,3709,4128,4952,4994,6589,8232,8250,9469,10674,12349,12629,14869,15229,
69,120,830,1479,3498,3710,4129,4953,4995,6590,8233,8251,9470,10675,12350,12630,14870,15230,
70,121,831,1480,3499,3711,4130,4954,4996,6591,8234,8252,9471,10676,12351,12631,14871,15231,
71,122,832,1481,3500,3712,4131,4955,4997,6592,8235,8253,9472,10677,12352,12632,14872,15232,
72,123,833,1482,3501,3713,4132,4956,4998,6593,8236,8254,9473,10678,12353,12633,14873,15233,
73,124,834,1483,3502,3714,4133,4957,4999,6594,8237,8255,9474,10679,12354,12634,14874,15234,
74,125,835,1484,3503,3715,4134,4958,5000,6595,8238,8256,9475,10680,12355,12635,14875,15235,
75,126,836,1485,3504,3716,4135,4959,5001,6596,8239,8257,9476,10681,12356,12636,14876,15236,
76,127,837,1486,3505,3717,4136,4960,5002,6597,8240,8258,9477,10682,12357,12637,14877,15237,
77,128,838,1487,3506,3718,4137,4961,5003,6598,8241,8259,9478,10683,12358,12638,14878,15238,
78,129,839,1488,3507,3719,4138,4962,5004,6599,8242,8260,9479,10684,12359,12639,14879,15239,
79,130,840,1489,3508,3720,4139,4963,5005,6600,8243,8261,9480,10685,12360,12640,14880,15240,
80,131,841,1490,3509,3721,4140,4964,5006,6601,8244,8262,9481,10686,12361,12641,14881,15241,
81,132,842,1491,3510,3722,4141,4965,5007,6602,8245,8263,9482,10687,12362,12642,14882,15242,
82,133,843,1492,3511,3723,4142,4966,5008,6603,8246,8264,9483,10688,12363,12643,14883,15243,
83,134,844,1493,3512,3724,4143,4967,5009,6604,8247,8265,9484,10689,12364,12644,14884,15244,
84,135,845,1494,3513,3725,4144,4968,5010,6605,8248,8266,9485,10690,12365,12645,14885,15245,
85,136,846,1495,3514,3726,4145,4969,5011,6606,8249,8267,9486,10691,12366,12646,14886,15246,
86,137,847,1496,3515,3727,4146,4970,5012,6607,8250,8268,9487,10692,12367,12647,14887,15247,
87,138,848,1497,3516,3728,4147,4971,5013,6608,8251,8269,9488,10693,12368,12648,14888,15248,
88,139,849,1498,3517,3729,4148,4972,5014,6609,8252,8270,9489,10694,12369,12649,14889,15249,
89,140,850,1499,3518,3730,4149,4973,5015,6610,8253,8271,9490,10695,12370,12650,14890,15250,
90,141,851,1500,3519,3731,4150,4974,5016,6611,8254,8272,9491,10696,12371,12651,14891,15251,
91,142,852,1501,3520,3732,4151,4975,5017,6612,8255,8273,9492,10697,12372,12652,14892,15252,
92,143,853,1502,3521,3733,4152,4976,5018,6613,8256,8274,9493,10698,12373,12653,14893,15253,
93,144,854,1503,3522,3734,4153,4977,5019,6614,8257,8275,9494,10699,12374,12654,14894,15254,
94,145,855,1504,3523,3735,4154,4978,5020,6615,8258,8276,9495,10700,12375,12655,14895,15255,
95,146,856,1505,3524,3736,4155,4979,5021,6616,8259,8277,9496,10701,12376,12656,14896,15256,
96,147,857,1506,3525,3737,4156,4980,5022,6617,8260,8278,9497,10702,12377,12657,14897,15257,
97,148,858,1507,3526,3738,4157,4981,5023,6618,8261,8279,9498,10703,12378,12658,14898,15258,
98,149,859,1508,3527,3739,4158,4982,5024,6619,7920,8262,9499,10704,12379,12659,14899,15259,
99,150,860,1509,3528,3740,4159,4983,5025,6620,7921,8263,9500,10705,12380,12660,14900,15260,
100,151,861,1510,3529,3741,4160,4984,5026,6621,7922,8264,9501,10706,12381,12661,14901,15261,
101,152,862,1511,3530,3742,4161,4985,5027,6622,7923,8265,9502,10707,12382,12662,14902,15262,
102,153,863,1512,3531,3743,4162,4986,5028,6623,7924,8266,9503,10708,12383,12663,14903,15263,
103,154,864,1513,3532,3744,4163,4987,5029,6624,7925,8267,9504,10709,12384,12664,14904,15264,
104,155,865,1514,3533,3745,4164,4988,5030,6625,7926,8268,9505,10710,12385,12665,14905,15265,
105,156,866,1515,3534,3746,4165,4989,5031,6626,7927,8269,9506,10711,12386,12666,14906,15266,
106,157,867,1516,3535,3747,4166,4990,5032,6627,7928,8270,9507,10712,12387,12667,14907,15267,
107,158,868,1517,3536,3748,4167,4991,5033,6628,7929,8271,9508,10713,12388,12668,14908,15268,
108,159,869,1518,3537,3749,4168,4992,5034,6629,7930,8272,9509,10714,12389,12669,14909,15269,
109,160,870,1519,3538,3750,4169,4993,5035,6630,7931,8273,9510,10715,12390,12670,14910,15270,
110,161,871,1520,3539,3751,4170,4994,5036,6631,7932,8274,9511,10716,12391,12671,14911,15271,
111,162,872,1521,3540,3752,4171,4995,5037,6632,7933,8275,9512,10717,12392,12672,14912,15272,
112,163,873,1522,3541,3753,4172,4996,5038,6633,7934,8276,9513,10718,12393,12673,14913,15273,
113,164,874,1523,3542,3754,4173,4997,5039,6634,7935,8277,9514,10719,12394,12674,14914,15274,
114,165,875,1524,3543,3755,4174,4680,4998,6635,7936,8278,9515,10720,12395,12675,14915,15275,
115,166,876,1525,3544,3756,4175,4681,4999,6636,7937,8279,9516,10721,12396,12676,14916,15276,
116,167,877,1526,3545,3757,4176,4682,5000,6637,7920,7938,9517,10722,12397,12677,14917,15277,
117,168,878,1527,3546,3758,4177,4683,5001,6638,7921,7939,9518,10723,12398,12678,14918,15278,
118,169,879,1528,3547,3759,4178,4684,5002,6639,7922,7940,9519,10724,12399,12679,14919,15279,
119,170,880,1529,3548,3760,4179,4685,5003,6640,7923,7941,9520,10725,12400,12680,14920,15280,
120,171,881,1530,3549,3761,4180,4686,5004,6641,7924,7942,9521,10726,12401,12681,14921,15281,
121,172,882,1531,3550,3762,4181,4687,5005,6642,7925,7943,9522,10727,12402,12682,14922,15282,
122,173,883,1532,3551,3763,4182,4688,5006,6643,7926,7944,9523,10728,12403,12683,14923,15283,
123,174,884,1533,3552,3764,4183,4689,5007,6644,7927,7945,9524,10729,12404,12684,14924,15284,
124,175,885,1534,3553,3765,4184,4690,5008,6645,7928,7946,9525,10730,12405,12685,14925,15285,
125,176,886,1535,3554,3766,4185,4691,5009,6646,7929,7947,9526,10731,12406,12686,14926,15286,
126,177,887,1536,3555,3767,4186,4692,5010,6647,7930,7948,9527,10732,12407,12687,14927,15287,
127,178,888,1537,3556,3768,4187,4693,5011,6648,7931,7949,9528,10733,12408,12688,14928,15288,
128,179,889,1538,3557,3769,4188,4694,5012,6649,7932,7950,9529,10734,12409,12689,14929,15289,
129,180,890,1539,3558,3770,4189,4695,5013,6650,7933,7951,9530,10735,12410,12690,14930,15290,
130,181,891,1540,3559,3771,4190,4696,5014,6651,7934,7952,9531,10736,12411,12691,14931,15291,
131,182,892,1541,3560,3772,4191,4697,5015,6652,7935,7953,9532,10737,12412,12692,14932,15292,
132,183,893,1542,3561,3773,4192,4698,5016,6653,7936,7954,9533,10738,12413,12693,14933,15293,
133,184,894,1543,3562,3774,4193,4699,5017,6654,7937,7955,9534,10739,12414,12694,14934,15294,
134,185,895,1544,3563,3775,4194,4700,5018,6655,7938,7956,9535,10740,12415,12695,14935,15295,
135,186,896,1545,3564,3776,4195,4701,5019,6656,7939,7957,9536,10741,12416,12696,14936,15296,
136,187,897,1546,3565,3777,4196,4702,5020,6657,7940,7958,9537,10742,12417,12697,14937,15297,
137,188,898,1547,3566,3778,4197,4703,5021,6658,7941,7959,9538,10743,12418,12698,14938,15298,
138,189,899,1548,3567,3779,4198,4704,5022,6659,7942,7960,9539,10744,12419,12699,14939,15299,
139,190,900,1549,3568,3780,4199,4705,5023,6660,7943,7961,9540,10745,12420,12700,14940,15300,
140,191,901,1550,3569,3781,4200,4706,5024,6661,7944,7962,9541,10746,12421,12701,14941,15301,
141,192,902,1551,3570,3782,4201,4707,5025,6662,7945,7963,9542,10747,12422,12702,14942,15302,
142,193,903,1552,3571,3783,4202,4708,5026,6663,7946,7964,9543,10748,12423,12703,14943,15303,
143,194,904,1553,3572,3784,4203,4709,5027,6664,7947,7965,9544,10749,12424,12704,14944,15304,
144,195,905,1554,3573,3785,4204,4710,5028,6665,7948,7966,9545,10750,12425,12705,14945,15305,
145,196,906,1555,3574,3786,4205,4711,5029,6666,7949,7967,9546,10751,12426,12706,14946,15306,
146,197,907,1556,3575,3787,4206,4712,5030,6667,7950,7968,9547,10752,12427,12707,14947,15307,
147,198,908,1557,3576,3788,4207,4713,5031,6668,7951,7969,9548,10753,12428,12708,14948,15308,
148,199,909,1558,3577,3789,4208,4714,5032,6669,7952,7970,9549,10754,12429,12709,14949,15309,
149,200,910,1559,3578,3790,4209,4715,5033,6670,7953,7971,9550,10755,12430,12710,14950,15310,
150,201,911,1560,3579,3791,4210,4716,5034,6671,7954,7972,9551,10756,12431,12711,14951,15311,
151,202,912,1561,3580,3792,4211,4717,5035,6672,7955,7973,9552,10757,12432,12712,14952,15312,
152,203,913,1562,3581,3793,4212,4718,5036,6673,7956,7974,9553,10758,12433,12713,14953,15313,
153,204,914,1563,3582,3794,4213,4719,5037,6674,7957,7975,9554,10759,12434,12714,14954,15314,
154,205,915,1564,3583,3795,4214,4720,5038,6675,7958,7976,9555,10760,12435,12715,14955,15315,
155,206,916,1565,3584,3796,4215,4721,5039,6676,7959,7977,9556,10761,12436,12716,14956,15316,
156,207,917,1566,3585,3797,4216,4680,4722,6677,7960,7978,9557,10762,12437,12717,14957,15317,
157,208,918,1567,3586,3798,4217,4681,4723,6678,7961,7979,9558,10763,12438,12718,14958,15318,
158,209,919,1568,3587,3799,4218,4682,4724,6679,7962,7980,9559,10764,12439,12719,14959,15319,
159,210,920,1569,3588,3800,4219,4683,4725,6680,7963,7981,9560,10765,12440,12720,14960,15320,
160,211,921,1570,3589,3801,4220,4684,4726,6681,7964,7982,9561,10766,12441,12721,14961,15321,
161,212,922,1571,3590,3802,4221,4685,4727,6682,7965,7983,9562,10767,12442,12722,14962,15322,
162,213,923,1572,3591,3803,4222,4686,4728,6683,7966,7984,9563,10768,12443,12723,14963,15323,
163,214,924,1573,3592,3804,4223,4687,4729,6684,7967,7985,9564,10769,12444,12724,14964,15324,
164,215,925,1574,3593,3805,4224,4688,4730,6685,7968,7986,9565,10770,12445,12725,14965,15325,
165,216,926,1575,3594,3806,4225,4689,4731,6686,7969,7987,9566,10771,12446,12726,14966,15326,
166,217,927,1576,3595,3807,4226,4690,4732,6687,7970,7988,9567,10772,12447,12727,14967,15327,
167,218,928,1577,3596,3808,4227,4691,4733,6688,7971,7989,9568,10773,12448,12728,14968,15328,
168,219,929,1578,3597,3809,4228,4692,4734,6689,7972,7990,9569,10774,12449,12729,14969,15329,
169,220,930,1579,3598,3810,4229,4693,4735,6690,7973,7991,9570,10775,12450,12730,14970,15330,
170,221,931,1580,3599,3811,4230,4694,4736,6691,7974,7992,9571,10776,12451,12731,14971,15331,
171,222,932,1581,3240,3812,4231,4695,4737,6692,7975,7993,9572,10777,12452,12732,14972,15332,
172,223,933,1582,3241,3813,4232,4696,4738,6693,7976,7994,9573,10778,12453,12733,14973,15333,
173,224,934,1583,3242,3814,4233,4697,4739,6694,7977,7995,9574,10779,12454,12734,14974,15334,
174,225,935,1584,3243,3815,4234,4698,4740,6695,7978,7996,9575,10780,12455,12735,14975,15335,
175,226,936,1585,3244,3816,4235,4699,4741,6696,7979,7997,9576,10781,12456,12736,14976,15336,
176,227,937,1586,3245,3817,4236,4700,4742,6697,7980,7998,9577,10782,12457,12737,14977,15337,
177,228,938,1587,3246,3818,4237,4701,4743,6698,7981,7999,9578,10783,12458,12738,14978,15338,
178,229,939,1588,3247,3819,4238,4702,4744,6699,7982,8000,9579,10784,12459,12739,14979,15339,
179,230,940,1589,3248,3820,4239,4703,4745,6700,7983,8001,9580,10785,12460,12740,14980,15340,
180,231,941,1590,3249,3821,4240,4704,4746,6701,7984,8002,9581,10786,12461,12741,14981,15341,
181,232,942,1591,3250,3822,4241,4705,4747,6702,7985,8003,9582,10787,12462,12742,14982,15342,
182,233,943,1592,3251,3823,4242,4706,4748,6703,7986,8004,9583,10788,12463,12743,14983,15343,
183,234,944,1593,3252,3824,4243,4707,4749,6704,7987,8005,9584,10789,12464,12744,14984,15344,
184,235,945,1594,3253,3825,4244,4708,4750,6705,7988,8006,9585,10790,12465,12745,14985,15345,
185,236,946,1595,3254,3826,4245,4709,4751,6706,7989,8007,9586,10791,12466,12746,14986,15346,
186,237,947,1596,3255,3827,4246,4710,4752,6707,7990,8008,9587,10792,12467,12747,14987,15347,
187,238,948,1597,3256,3828,4247,4711,4753,6708,7991,8009,9588,10793,12468,12748,14988,15348,
188,239,949,1598,3257,3829,4248,4712,4754,6709,7992,8010,9589,10794,12469,12749,14989,15349,
189,240,950,1599,3258,3830,4249,4713,4755,6710,7993,8011,9590,10795,12470,12750,14990,15350,
190,241,951,1600,3259,3831,4250,4714,4756,6711,7994,8012,9591,10796,12471,12751,14991,15351,
191,242,952,1601,3260,3832,4251,4715,4757,6712,7995,8013,9592,10797,12472,12752,14992,15352,
192,243,953,1602,3261,3833,4252,4716,4758,6713,7996,8014,9593,10798,12473,12753,14993,15353,
193,244,954,1603,3262,3834,4253,4717,4759,6714,7997,8015,9594,10799,12474,12754,14994,15354,
194,245,955,1604,3263,3835,4254,4718,4760,6715,7998,8016,9595,10440,12475,12755,14995,15355,
195,246,956,1605,3264,3836,4255,4719,4761,6716,7999,8017,9596,10441,12476,12756,14996,15356,
196,247,957,1606,3265,3837,4256,4720,4762,6717,8000,8018,9597,10442,12477,12757,14997,15357,
197,248,958,1607,3266,3838,4257,4721,4763,6718,8001,8019,9598,10443,12478,12758,14998,15358,
198,249,959,1608,3267,3839,4258,4722,4764,6719,8002,8020,9599,10444,12479,12759,14999,15359,
199,250,960,1609,3268,3840,4259,4723,4765,6720,8003,8021,9600,10445,12480,12760,15000,15360,
200,251,961,1610,3269,3841,4260,4724,4766,6721,8004,8022,9601,10446,12481,12761,15001,15361,
201,252,962,1611,3270,3842,4261,4725,4767,6722,8005,8023,9602,10447,12482,12762,15002,15362,
202,253,963,1612,3271,3843,4262,4726,4768,6723,8006,8024,9603,10448,12483,12763,15003,15363,
203,254,964,1613,3272,3844,4263,4727,4769,6724,8007,8025,9604,10449,12484,12764,15004,15364,
204,255,965,1614,3273,3845,4264,4728,4770,6725,8008,8026,9605,10450,12485,12765,15005,15365,
205,256,966,1615,3274,3846,4265,4729,4771,6726,8009,8027,9606,10451,12486,12766,15006,15366,
206,257,967,1616,3275,3847,4266,4730,4772,6727,8010,8028,9607,10452,12487,12767,15007,15367,
207,258,968,1617,3276,3848,4267,4731,4773,6728,8011,8029,9608,10453,12488,12768,15008,15368,
208,259,969,1618,3277,3849,4268,4732,4774,6729,8012,8030,9609,10454,12489,12769,15009,15369,
209,260,970,1619,3278,3850,4269,4733,4775,6730,8013,8031,9610,10455,12490,12770,15010,15370,
210,261,971,1620,3279,3851,4270,4734,4776,6731,8014,8032,9611,10456,12491,12771,15011,15371,
211,262,972,1621,3280,3852,4271,4735,4777,6732,8015,8033,9612,10457,12492,12772,15012,15372,
212,263,973,1622,3281,3853,4272,4736,4778,6733,8016,8034,9613,10458,12493,12773,15013,15373,
213,264,974,1623,3282,3854,4273,4737,4779,6734,8017,8035,9614,10459,12494,12774,15014,15374,
214,265,975,1624,3283,3855,4274,4738,4780,6735,8018,8036,9615,10460,12495,12775,15015,15375,
215,266,976,1625,3284,3856,4275,4739,4781,6736,8019,8037,9616,10461,12496,12776,15016,15376,
216,267,977,1626,3285,3857,4276,4740,4782,6737,8020,8038,9617,10462,12497,12777,15017,15377,
217,268,978,1627,3286,3858,4277,4741,4783,6738,8021,8039,9618,10463,12498,12778,15018,15378,
218,269,979,1628,3287,3859,4278,4742,4784,6739,8022,8040,9619,10464,12499,12779,15019,15379,
219,270,980,1629,3288,3860,4279,4743,4785,6740,8023,8041,9620,10465,12500,12780,15020,15380,
220,271,981,1630,3289,3861,4280,4744,4786,6741,8024,8042,9621,10466,12501,12781,15021,15381,
221,272,982,1631,3290,3862,4281,4745,4787,6742,8025,8043,9622,10467,12502,12782,15022,15382,
222,273,983,1632,3291,3863,4282,4746,4788,6743,8026,8044,9623,10468,12503,12783,15023,15383,
223,274,984,1633,3292,3864,4283,4747,4789,6744,8027,8045,9624,10469,12504,12784,15024,15384,
224,275,985,1634,3293,3865,4284,4748,4790,6745,8028,8046,9625,10470,12505,12785,15025,15385,
225,276,986,1635,3294,3866,4285,4749,4791,6746,8029,8047,9626,10471,12506,12786,15026,15386,
226,277,987,1636,3295,3867,4286,4750,4792,6747,8030,8048,9627,10472,12507,12787,15027,15387,
227,278,988,1637,3296,3868,4287,4751,4793,6748,8031,8049,9628,10473,12508,12788,15028,15388,
228,279,989,1638,3297,3869,4288,4752,4794,6749,8032,8050,9629,10474,12509,12789,15029,15389,
229,280,990,1639,3298,3870,4289,4753,4795,6750,8033,8051,9630,10475,12510,12790,15030,15390,
230,281,991,1640,3299,3871,4290,4754,4796,6751,8034,8052,9631,10476,12511,12791,15031,15391,
231,282,992,1641,3300,3872,4291,4755,4797,6752,8035,8053,9632,10477,12512,12792,15032,15392,
232,283,993,1642,3301,3873,4292,4756,4798,6753,8036,8054,9633,10478,12513,12793,15033,15393,
233,284,994,1643,3302,3874,4293,4757,4799,6754,8037,8055,9634,10479,12514,12794,15034,15394,
234,285,995,1644,3303,3875,4294,4758,4800,6755,8038,8056,9635,10480,12515,12795,15035,15395,
235,286,996,1645,3304,3876,4295,4759,4801,6756,8039,8057,9636,10481,12516,12796,15036,15396,
236,287,997,1646,3305,3877,4296,4760,4802,6757,8040,8058,9637,10482,12517,12797,15037,15397,
237,288,998,1647,3306,3878,4297,4761,4803,6758,8041,8059,9638,10483,12518,12798,15038,15398,
238,289,999,1648,3307,3879,4298,4762,4804,6759,8042,8060,9639,10484,12519,12799,15039,15399,
239,290,1000,1649,3308,3880,4299,4763,4805,6760,8043,8061,9640,10485,12520,12800,15040,15400,
240,291,1001,1650,3309,3881,4300,4764,4806,6761,8044,8062,9641,10486,12521,12801,15041,15401,
241,292,1002,1651,3310,3882,4301,4765,4807,6762,8045,8063,9642,10487,12522,12802,15042,15402,
242,293,1003,1652,3311,3883,4302,4766,4808,6763,8046,8064,9643,10488,12523,12803,15043,15403,
243,294,1004,1653,3312,3884,4303,4767,4809,6764,8047,8065,9644,10489,12524,12804,15044,15404,
244,295,1005,1654,3313,3885,4304,4768,4810,6765,8048,8066,9645,10490,12525,12805,15045,15405,
245,296,1006,1655,3314,3886,4305,4769,4811,6766,8049,8067,9646,10491,12526,12806,15046,15406,
246,297,1007,1656,3315,3887,4306,4770,4812,6767,8050,8068,9647,10492,12527,12807,15047,15407,
247,298,1008,1657,3316,3888,4307,4771,4813,6768,8051,8069,9648,10493,12528,12808,15048,15408,
248,299,1009,1658,3317,3889,4308,4772,4814,6769,8052,8070,9649,10494,12529,12809,15049,15409,
249,300,1010,1659,3318,3890,4309,4773,4815,6770,8053,8071,9650,10495,12530,12810,15050,15410,
250,301,1011,1660,3319,3891,4310,4774,4816,6771,8054,8072,9651,10496,12531,12811,15051,15411,
251,302,1012,1661,3320,3892,4311,4775,4817,6772,8055,8073,9652,10497,12532,12812,15052,15412,
252,303,1013,1662,3321,3893,4312,4776,4818,6773,8056,8074,9653,10498,12533,12813,15053,15413,
253,304,1014,1663,3322,3894,4313,4777,4819,6774,8057,8075,9654,10499,12534,12814,15054,15414,
254,305,1015,1664,3323,3895,4314,4778,4820,6775,8058,8076,9655,10500,12535,12815,15055,15415,
255,306,1016,1665,3324,3896,4315,4779,4821,6776,8059,8077,9656,10501,12536,12816,15056,15416,
256,307,1017,1666,3325,3897,4316,4780,4822,6777,8060,8078,9657,10502,12537,12817,15057,15417,
257,308,1018,1667,3326,3898,4317,4781,4823,6778,8061,8079,9658,10503,12538,12818,15058,15418,
258,309,1019,1668,3327,3899,4318,4782,4824,6779,8062,8080,9659,10504,12539,12819,15059,15419,
259,310,1020,1669,3328,3900,4319,4783,4825,6780,8063,8081,9660,10505,12540,12820,15060,15420,
260,311,1021,1670,3329,3901,3960,4784,4826,6781,8064,8082,9661,10506,12541,12821,15061,15421,
261,312,1022,1671,3330,3902,3961,4785,4827,6782,8065,8083,9662,10507,12542,12822,15062,15422,
262,313,1023,1672,3331,3903,3962,4786,4828,6783,8066,8084,9663,10508,12543,12823,15063,15423,
263,314,1024,1673,3332,3904,3963,4787,4829,6784,8067,8085,9664,10509,12544,12824,15064,15424,
264,315,1025,1674,3333,3905,3964,4788,4830,6785,8068,8086,9665,10510,12545,12825,15065,15425,
265,316,1026,1675,3334,3906,3965,4789,4831,6786,8069,8087,9666,10511,12546,12826,15066,15426,
266,317,1027,1676,3335,3907,3966,4790,4832,6787,8070,8088,9667,10512,12547,12827,15067,15427,
267,318,1028,1677,3336,3908,3967,4791,4833,6788,8071,8089,9668,10513,12548,12828,15068,15428,
268,319,1029,1678,3337,3909,3968,4792,4834,6789,8072,8090,9669,10514,12549,12829,15069,15429,
269,320,1030,1679,3338,3910,3969,4793,4835,6790,8073,8091,9670,10515,12550,12830,15070,15430,
270,321,1031,1680,3339,3911,3970,4794,4836,6791,8074,8092,9671,10516,12551,12831,15071,15431,
271,322,1032,1681,3340,3912,3971,4795,4837,6792,8075,8093,9672,10517,12552,12832,15072,15432,
272,323,1033,1682,3341,3913,3972,4796,4838,6793,8076,8094,9673,10518,12553,12833,15073,15433,
273,324,1034,1683,3342,3914,3973,4797,4839,6794,8077,8095,9674,10519,12554,12834,15074,15434,
274,325,1035,1684,3343,3915,3974,4798,4840,6795,8078,8096,9675,10520,12555,12835,15075,15435,
275,326,1036,1685,3344,3916,3975,4799,4841,6796,8079,8097,9676,10521,12556,12836,15076,15436,
276,327,1037,1686,3345,3917,3976,4800,4842,6797,8080,8098,9677,10522,12557,12837,15077,15437,
277,328,1038,1687,3346,3918,3977,4801,4843,6798,8081,8099,9678,10523,12558,12838,15078,15438,
278,329,1039,1688,3347,3919,3978,4802,4844,6799,8082,8100,9679,10524,12559,12839,15079,15439,
279,330,1040,1689,3348,3920,3979,4803,4845,6800,8083,8101,9680,10525,12560,12840,15080,15440,
280,331,1041,1690,3349,3921,3980,4804,4846,6801,8084,8102,9681,10526,12561,12841,15081,15441,
281,332,1042,1691,3350,3922,3981,4805,4847,6802,8085,8103,9682,10527,12562,12842,15082,15442,
282,333,1043,1692,3351,3923,3982,4806,4848,6803,8086,8104,9683,10528,12563,12843,15083,15443,
283,334,1044,1693,3352,3924,3983,4807,4849,6804,8087,8105,9684,10529,12564,12844,15084,15444,
284,335,1045,1694,3353,3925,3984,4808,4850,6805,8088,8106,9685,10530,12565,12845,15085,15445,
285,336,1046,1695,3354,3926,3985,4809,4851,6806,8089,8107,9686,10531,12566,12846,15086,15446,
286,337,1047,1696,3355,3927,3986,4810,4852,6807,8090,8108,9687,10532,12567,12847,15087,15447,
287,338,1048,1697,3356,3928,3987,4811,4853,6808,8091,8109,9688,10533,12568,12848,15088,15448,
288,339,1049,1698,3357,3929,3988,4812,4854,6809,8092,8110,9689,10534,12569,12849,15089,15449,
289,340,1050,1699,3358,3930,3989,4813,4855,6810,8093,8111,9690,10535,12570,12850,15090,15450,
290,341,1051,1700,3359,3931,3990,4814,4856,6811,8094,8112,9691,10536,12571,12851,15091,15451,
291,342,1052,1701,3360,3932,3991,4815,4857,6812,8095,8113,9692,10537,12572,12852,15092,15452,
292,343,1053,1702,3361,3933,3992,4816,4858,6813,8096,8114,9693,10538,12573,12853,15093,15453,
293,344,1054,1703,3362,3934,3993,4817,4859,6814,8097,8115,9694,10539,12574,12854,15094,15454,
294,345,1055,1704,3363,3935,3994,4818,4860,6815,8098,8116,9695,10540,12575,12855,15095,15455,
295,346,1056,1705,3364,3936,3995,4819,4861,6816,8099,8117,9696,10541,12576,12856,15096,15456,
296,347,1057,1706,3365,3937,3996,4820,4862,6817,8100,8118,9697,10542,12577,12857,15097,15457,
297,348,1058,1707,3366,3938,3997,4821,4863,6818,8101,8119,9698,10543,12578,12858,15098,15458,
298,349,1059,1708,3367,3939,3998,4822,4864,6819,8102,8120,9699,10544,12579,12859,15099,15459,
299,350,1060,1709,3368,3940,3999,4823,4865,6820,8103,8121,9700,10545,12580,12860,15100,15460,
300,351,1061,1710,3369,3941,4000,4824,4866,6821,8104,8122,9701,10546,12581,12861,15101,15461,
301,352,1062,1711,3370,3942,4001,4825,4867,6822,8105,8123,9702,10547,12582,12862,15102,15462,
302,353,1063,1712,3371,3943,4002,4826,4868,6823,8106,8124,9703,10548,12583,12863,15103,15463,
303,354,1064,1713,3372,3944,4003,4827,4869,6824,8107,8125,9704,10549,12584,12864,15104,15464,
304,355,1065,1714,3373,3945,4004,4828,4870,6825,8108,8126,9705,10550,12585,12865,15105,15465,
305,356,1066,1715,3374,3946,4005,4829,4871,6826,8109,8127,9706,10551,12586,12866,15106,15466,
306,357,1067,1716,3375,3947,4006,4830,4872,6827,8110,8128,9707,10552,12587,12867,15107,15467,
307,358,1068,1717,3376,3948,4007,4831,4873,6828,8111,8129,9708,10553,12588,12868,15108,15468,
308,359,1069,1718,3377,3949,4008,4832,4874,6829,8112,8130,9709,10554,12589,12869,15109,15469,
0,309,1070,1719,3378,3950,4009,4833,4875,6830,8113,8131,9710,10555,12590,12870,15110,15470,
1,310,1071,1720,3379,3951,4010,4834,4876,6831,8114,8132,9711,10556,12591,12871,15111,15471,
2,311,1072,1721,3380,3952,4011,4835,4877,6832,8115,8133,9712,10557,12592,12872,15112,15472,
3,312,1073,1722,3381,3953,4012,4836,4878,6833,8116,8134,9713,10558,12593,12873,15113,15473,
4,313,1074,1723,3382,3954,4013,4837,4879,6834,8117,8135,9714,10559,12594,12874,15114,15474,
5,314,1075,1724,3383,3955,4014,4838,4880,6835,8118,8136,9715,10560,12595,12875,15115,15475,
6,315,1076,1725,3384,3956,4015,4839,4881,6836,8119,8137,9716,10561,12596,12876,15116,15476,
7,316,1077,1726,3385,3957,4016,4840,4882,6837,8120,8138,9717,10562,12597,12877,15117,15477,
8,317,1078,1727,3386,3958,4017,4841,4883,6838,8121,8139,9718,10563,12598,12878,15118,15478,
9,318,1079,1728,3387,3959,4018,4842,4884,6839,8122,8140,9719,10564,12599,12879,15119,15479,
148,202,480,1029,1080,2235,3940,3960,6719,6840,7270,8816,9720,9921,11416,11632,12600,15120,15480,
149,203,481,1030,1081,2236,3941,3961,6720,6841,7271,8817,9721,9922,11417,11633,12601,15121,15481,
150,204,482,1031,1082,2237,3942,3962,6721,6842,7272,8818,9722,9923,11418,11634,12602,15122,15482,
151,205,483,1032,1083,2238,3943,3963,6722,6843,7273,8819,9723,9924,11419,11635,12603,15123,15483,
152,206,484,1033,1084,2239,3944,3964,6723,6844,7274,8820,9724,9925,11420,11636,12604,15124,15484,
153,207,485,1034,1085,2240,3945,3965,6724,6845,7275,8821,9725,9926,11421,11637,12605,15125,15485,
154,208,486,1035,1086,2241,3946,3966,6725,6846,7276,8822,9726,9927,11422,11638,12606,15126,15486,
155,209,487,1036,1087,2242,3947,3967,6726,6847,7277,8823,9727,9928,11423,11639,12607,15127,15487,
156,210,488,1037,1088,2243,3948,3968,6727,6848,7278,8824,9728,9929,11424,11640,12608,15128,15488,
157,211,489,1038,1089,2244,3949,3969,6728,6849,7279,8825,9729,9930,11425,11641,12609,15129,15489,
158,212,490,1039,1090,2245,3950,3970,6729,6850,7280,8826,9730,9931,11426,11642,12610,15130,15490,
159,213,491,1040,1091,2246,3951,3971,6730,6851,7281,8827,9731,9932,11427,11643,12611,15131,15491,
160,214,492,1041,1092,2247,3952,3972,6731,6852,7282,8828,9732,9933,11428,11644,12612,15132,15492,
161,215,493,1042,1093,2248,3953,3973,6732,6853,7283,8829,9733,9934,11429,11645,12613,15133,15493,
162,216,494,1043,1094,2249,3954,3974,6733,6854,7284,8830,9734,9935,11430,11646,12614,15134,15494,
163,217,495,1044,1095,2250,3955,3975,6734,6855,7285,8831,9735,9936,11431,11647,12615,15135,15495,
164,218,496,1045,1096,2251,3956,3976,6735,6856,7286,8832,9736,9937,11432,11648,12616,15136,15496,
165,219,497,1046,1097,2252,3957,3977,6736,6857,7287,8833,9737,9938,11433,11649,12617,15137,15497,
166,220,498,1047,1098,2253,3958,3978,6737,6858,7288,8834,9738,9939,11434,11650,12618,15138,15498,
167,221,499,1048,1099,2254,3959,3979,6738,6859,7289,8835,9739,9940,11435,11651,12619,15139,15499,
168,222,500,1049,1100,2255,3600,3980,6739,6860,7290,8836,9740,9941,11436,11652,12620,15140,15500,
169,223,501,1050,1101,2256,3601,3981,6740,6861,7291,8837,9741,9942,11437,11653,12621,15141,15501,
170,224,502,1051,1102,2257,3602,3982,6741,6862,7292,8838,9742,9943,11438,11654,12622,15142,15502,
171,225,503,1052,1103,2258,3603,3983,6742,6863,7293,8839,9743,9944,11439,11655,12623,15143,15503,
172,226,504,1053,1104,2259,3604,3984,6743,6864,7294,8840,9744,9945,11440,11656,12624,15144,15504,
173,227,505,1054,1105,2260,3605,3985,6744,6865,7295,8841,9745,9946,11441,11657,12625,15145,15505,
174,228,506,1055,1106,2261,3606,3986,6745,6866,7296,8842,9746,9947,11442,11658,12626,15146,15506,
175,229,507,1056,1107,2262,3607,3987,6746,6867,7297,8843,9747,9948,11443,11659,12627,15147,15507,
176,230,508,1057,1108,2263,3608,3988,6747,6868,7298,8844,9748,9949,11444,11660,12628,15148,15508,
177,231,509,1058,1109,2264,3609,3989,6748,6869,7299,8845,9749,9950,11445,11661,12629,15149,15509,
178,232,510,1059,1110,2265,3610,3990,6749,6870,7300,8846,9750,9951,11446,11662,12630,15150,15510,
179,233,511,1060,1111,2266,3611,3991,6750,6871,7301,8847,9751,9952,11447,11663,12631,15151,15511,
180,234,512,1061,1112,2267,3612,3992,6751,6872,7302,8848,9752,9953,11448,11664,12632,15152,15512,
181,235,513,1062,1113,2268,3613,3993,6752,6873,7303,8849,9753,9954,11449,11665,12633,15153,15513,
182,236,514,1063,1114,2269,3614,3994,6753,6874,7304,8850,9754,9955,11450,11666,12634,15154,15514,
183,237,515,1064,1115,2270,3615,3995,6754,6875,7305,8851,9755,9956,11451,11667,12635,15155,15515,
184,238,516,1065,1116,2271,3616,3996,6755,6876,7306,8852,9756,9957,11452,11668,12636,15156,15516,
185,239,517,1066,1117,2272,3617,3997,6756,6877,7307,8853,9757,9958,11453,11669,12637,15157,15517,
186,240,518,1067,1118,2273,3618,3998,6757,6878,7308,8854,9758,9959,11454,11670,12638,15158,15518,
187,241,519,1068,1119,2274,3619,3999,6758,6879,7309,8855,9759,9960,11455,11671,12639,15159,15519,
188,242,520,1069,1120,2275,3620,4000,6759,6880,7310,8856,9760,9961,11456,11672,12640,15160,15520,
189,243,521,1070,1121,2276,3621,4001,6760,6881,7311,8857,9761,9962,11457,11673,12641,15161,15521,
190,244,522,1071,1122,2277,3622,4002,6761,6882,7312,8858,9762,9963,11458,11674,12642,15162,15522,
191,245,523,1072,1123,2278,3623,4003,6762,6883,7313,8859,9763,9964,11459,11675,12643,15163,15523,
192,246,524,1073,1124,2279,3624,4004,6763,6884,7314,8860,9764,9965,11460,11676,12644,15164,15524,
193,247,525,1074,1125,2280,3625,4005,6764,6885,7315,8861,9765,9966,11461,11677,12645,15165,15525,
194,248,526,1075,1126,2281,3626,4006,6765,6886,7316,8862,9766,9967,11462,11678,12646,15166,15526,
195,249,527,1076,1127,2282,3627,4007,6766,6887,7317,8863,9767,9968,11463,11679,12647,15167,15527,
196,250,528,1077,1128,2283,3628,4008,6767,6888,7318,8864,9768,9969,11464,11680,12648,15168,15528,
197,251,529,1078,1129,2284,3629,4009,6768,6889,7319,8865,9769,9970,11465,11681,12649,15169,15529,
198,252,530,1079,1130,2285,3630,4010,6769,6890,7320,8866,9770,9971,11466,11682,12650,15170,15530,
199,253,531,720,1131,2286,3631,4011,6770,6891,7321,8867,9771,9972,11467,11683,12651,15171,15531,
200,254,532,721,1132,2287,3632,4012,6771,6892,7322,8868,9772,9973,11468,11684,12652,15172,15532,
201,255,533,722,1133,2288,3633,4013,6772,6893,7323,8869,9773,9974,11469,11685,12653,15173,15533,
202,256,534,723,1134,2289,3634,4014,6773,6894,7324,8870,9774,9975,11470,11686,12654,15174,15534,
203,257,535,724,1135,2290,3635,4015,6774,6895,7325,8871,9775,9976,11471,11687,12655,15175,15535,
204,258,536,725,1136,2291,3636,4016,6775,6896,7326,8872,9776,9977,11472,11688,12656,15176,15536,
205,259,537,726,1137,2292,3637,4017,6776,6897,7327,8873,9777,9978,11473,11689,12657,15177,15537,
206,260,538,727,1138,2293,3638,4018,6777,6898,7328,8874,9778,9979,11474,11690,12658,15178,15538,
207,261,539,728,1139,2294,3639,4019,6778,6899,7329,8875,9779,9980,11475,11691,12659,15179,15539,
208,262,540,729,1140,2295,3640,4020,6779,6900,7330,8876,9780,9981,11476,11692,12660,15180,15540,
209,263,541,730,1141,2296,3641,4021,6780,6901,7331,8877,9781,9982,11477,11693,12661,15181,15541,
210,264,542,731,1142,2297,3642,4022,6781,6902,7332,8878,9782,9983,11478,11694,12662,15182,15542,
211,265,543,732,1143,2298,3643,4023,6782,6903,7333,8879,9783,9984,11479,11695,12663,15183,15543,
212,266,544,733,1144,2299,3644,4024,6783,6904,7334,8880,9784,9985,11480,11696,12664,15184,15544,
213,267,545,734,1145,2300,3645,4025,6784,6905,7335,8881,9785,9986,11481,11697,12665,15185,15545,
214,268,546,735,1146,2301,3646,4026,6785,6906,7336,8882,9786,9987,11482,11698,12666,15186,15546,
215,269,547,736,1147,2302,3647,4027,6786,6907,7337,8883,9787,9988,11483,11699,12667,15187,15547,
216,270,548,737,1148,2303,3648,4028,6787,6908,7338,8884,9788,9989,11484,11700,12668,15188,15548,
217,271,549,738,1149,2304,3649,4029,6788,6909,7339,8885,9789,9990,11485,11701,12669,15189,15549,
218,272,550,739,1150,2305,3650,4030,6789,6910,7340,8886,9790,9991,11486,11702,12670,15190,15550,
219,273,551,740,1151,2306,3651,4031,6790,6911,7341,8887,9791,9992,11487,11703,12671,15191,15551,
220,274,552,741,1152,2307,3652,4032,6791,6912,7342,8888,9792,9993,11488,11704,12672,15192,15552,
221,275,553,742,1153,2308,3653,4033,6792,6913,7343,8889,9793,9994,11489,11705,12673,15193,15553,
222,276,554,743,1154,2309,3654,4034,6793,6914,7344,8890,9794,9995,11490,11706,12674,15194,15554,
223,277,555,744,1155,2310,3655,4035,6794,6915,7345,8891,9795,9996,11491,11707,12675,15195,15555,
224,278,556,745,1156,2311,3656,4036,6795,6916,7346,8892,9796,9997,11492,11708,12676,15196,15556,
225,279,557,746,1157,2312,3657,4037,6796,6917,7347,8893,9797,9998,11493,11709,12677,15197,15557,
226,280,558,747,1158,2313,3658,4038,6797,6918,7348,8894,9798,9999,11494,11710,12678,15198,15558,
227,281,559,748,1159,2314,3659,4039,6798,6919,7349,8895,9799,10000,11495,11711,12679,15199,15559,
228,282,560,749,1160,2315,3660,4040,6799,6920,7350,8896,9800,10001,11496,11712,12680,15200,15560,
229,283,561,750,1161,2316,3661,4041,6800,6921,7351,8897,9801,10002,11497,11713,12681,15201,15561,
230,284,562,751,1162,2317,3662,4042,6801,6922,7352,8898,9802,10003,11498,11714,12682,15202,15562,
231,285,563,752,1163,2318,3663,4043,6802,6923,7353,8899,9803,10004,11499,11715,12683,15203,15563,
232,286,564,753,1164,2319,3664,4044,6803,6924,7354,8900,9804,10005,11500,11716,12684,15204,15564,
233,287,565,754,1165,2320,3665,4045,6804,6925,7355,8901,9805,10006,11501,11717,12685,15205,15565,
234,288,566,755,1166,2321,3666,4046,6805,6926,7356,8902,9806,10007,11502,11718,12686,15206,15566,
235,289,567,756,1167,2322,3667,4047,6806,6927,7357,8903,9807,10008,11503,11719,12687,15207,15567,
236,290,568,757,1168,2323,3668,4048,6807,6928,7358,8904,9808,10009,11504,11720,12688,15208,15568,
237,291,569,758,1169,2324,3669,4049,6808,6929,7359,8905,9809,10010,11505,11721,12689,15209,15569,
238,292,570,759,1170,2325,3670,4050,6809,6930,7360,8906,9810,10011,11506,11722,12690,15210,15570,
239,293,571,760,1171,2326,3671,4051,6810,6931,7361,8907,9811,10012,11507,11723,12691,15211,15571,
240,294,572,761,1172,2327,3672,4052,6811,6932,7362,8908,9812,10013,11508,11724,12692,15212,15572,
241,295,573,762,1173,2328,3673,4053,6812,6933,7363,8909,9813,10014,11509,11725,12693,15213,15573,
242,296,574,763,1174,2329,3674,4054,6813,6934,7364,8910,9814,10015,11510,11726,12694,15214,15574,
243,297,575,764,1175,2330,3675,4055,6814,6935,7365,8911,9815,10016,11511,11727,12695,15215,15575,
244,298,576,765,1176,2331,3676,4056,6815,6936,7366,8912,9816,10017,11512,11728,12696,15216,15576,
245,299,577,766,1177,2332,3677,4057,6816,6937,7367,8913,9817,10018,11513,11729,12697,15217,15577,
246,300,578,767,1178,2333,3678,4058,6817,6938,7368,8914,9818,10019,11514,11730,12698,15218,15578,
247,301,579,768,1179,2334,3679,4059,6818,6939,7369,8915,9819,10020,11515,11731,12699,15219,15579,
248,302,580,769,1180,2335,3680,4060,6819,6940,7370,8916,9820,10021,11516,11732,12700,15220,15580,
249,303,581,770,1181,2336,3681,4061,6820,6941,7371,8917,9821,10022,11517,11733,12701,15221,15581,
250,304,582,771,1182,2337,3682,4062,6821,6942,7372,8918,9822,10023,11518,11734,12702,15222,15582,
251,305,583,772,1183,2338,3683,4063,6822,6943,7373,8919,9823,10024,11519,11735,12703,15223,15583,
252,306,584,773,1184,2339,3684,4064,6823,6944,7374,8920,9824,10025,11160,11736,12704,15224,15584,
253,307,585,774,1185,2340,3685,4065,6824,6945,7375,8921,9825,10026,11161,11737,12705,15225,15585,
254,308,586,775,1186,2341,3686,4066,6825,6946,7376,8922,9826,10027,11162,11738,12706,15226,15586,
255,309,587,776,1187,2342,3687,4067,6826,6947,7377,8923,9827,10028,11163,11739,12707,15227,15587,
256,310,588,777,1188,2343,3688,4068,6827,6948,7378,8924,9828,10029,11164,11740,12708,15228,15588,
257,311,589,778,1189,2344,3689,4069,6828,6949,7379,8925,9829,10030,11165,11741,12709,15229,15589,
258,312,590,779,1190,2345,3690,4070,6829,6950,7380,8926,9830,10031,11166,11742,12710,15230,15590,
259,313,591,780,1191,2346,3691,4071,6830,6951,7381,8927,9831,10032,11167,11743,12711,15231,15591,
260,314,592,781,1192,2347,3692,4072,6831,6952,7382,8928,9832,10033,11168,11744,12712,15232,15592,
261,315,593,782,1193,2348,3693,4073,6832,6953,7383,8929,9833,10034,11169,11745,12713,15233,15593,
262,316,594,783,1194,2349,3694,4074,6833,6954,7384,8930,9834,10035,11170,11746,12714,15234,15594,
263,317,595,784,1195,2350,3695,4075,6834,6955,7385,8931,9835,10036,11171,11747,12715,15235,15595,
264,318,596,785,1196,2351,3696,4076,6835,6956,7386,8932,9836,10037,11172,11748,12716,15236,15596,
265,319,597,786,1197,2352,3697,4077,6836,6957,7387,8933,9837,10038,11173,11749,12717,15237,15597,
266,320,598,787,1198,2353,3698,4078,6837,6958,7388,8934,9838,10039,11174,11750,12718,15238,15598,
267,321,599,788,1199,2354,3699,4079,6838,6959,7389,8935,9839,10040,11175,11751,12719,15239,15599,
268,322,600,789,1200,2355,3700,4080,6839,6960,7390,8936,9840,10041,11176,11752,12720,15240,15600,
269,323,601,790,1201,2356,3701,4081,6480,6961,7391,8937,9841,10042,11177,11753,12721,15241,15601,
270,324,602,791,1202,2357,3702,4082,6481,6962,7392,8938,9842,10043,11178,11754,12722,15242,15602,
271,325,603,792,1203,2358,3703,4083,6482,6963,7393,8939,9843,10044,11179,11755,12723,15243,15603,
272,326,604,793,1204,2359,3704,4084,6483,6964,7394,8940,9844,10045,11180,11756,12724,15244,15604,
273,327,605,794,1205,2360,3705,4085,6484,6965,7395,8941,9845,10046,11181,11757,12725,15245,15605,
274,328,606,795,1206,2361,3706,4086,6485,6966,7396,8942,9846,10047,11182,11758,12726,15246,15606,
275,329,607,796,1207,2362,3707,4087,6486,6967,7397,8943,9847,10048,11183,11759,12727,15247,15607,
276,330,608,797,1208,2363,3708,4088,6487,6968,7398,8944,9848,10049,11184,11760,12728,15248,15608,
277,331,609,798,1209,2364,3709,4089,6488,6969,7399,8945,9849,10050,11185,11761,12729,15249,15609,
278,332,610,799,1210,2365,3710,4090,6489,6970,7400,8946,9850,10051,11186,11762,12730,15250,15610,
279,333,611,800,1211,2366,3711,4091,6490,6971,7401,8947,9851,10052,11187,11763,12731,15251,15611,
280,334,612,801,1212,2367,3712,4092,6491,6972,7402,8948,9852,10053,11188,11764,12732,15252,15612,
281,335,613,802,1213,2368,3713,4093,6492,6973,7403,8949,9853,10054,11189,11765,12733,15253,15613,
282,336,614,803,1214,2369,3714,4094,6493,6974,7404,8950,9854,10055,11190,11766,12734,15254,15614,
283,337,615,804,1215,2370,3715,4095,6494,6975,7405,8951,9855,10056,11191,11767,12735,15255,15615,
284,338,616,805,1216,2371,3716,4096,6495,6976,7406,8952,9856,10057,11192,11768,12736,15256,15616,
285,339,617,806,1217,2372,3717,4097,6496,6977,7407,8953,9857,10058,11193,11769,12737,15257,15617,
286,340,618,807,1218,2373,3718,4098,6497,6978,7408,8954,9858,10059,11194,11770,12738,15258,15618,
287,341,619,808,1219,2374,3719,4099,6498,6979,7409,8955,9859,10060,11195,11771,12739,15259,15619,
288,342,620,809,1220,2375,3720,4100,6499,6980,7410,8956,9860,10061,11196,11772,12740,15260,15620,
289,343,621,810,1221,2376,3721,4101,6500,6981,7411,8957,9861,10062,11197,11773,12741,15261,15621,
290,344,622,811,1222,2377,3722,4102,6501,6982,7412,8958,9862,10063,11198,11774,12742,15262,15622,
291,345,623,812,1223,2378,3723,4103,6502,6983,7413,8959,9863,10064,11199,11775,12743,15263,15623,
292,346,624,813,1224,2379,3724,4104,6503,6984,7414,8960,9864,10065,11200,11776,12744,15264,15624,
293,347,625,814,1225,2380,3725,4105,6504,6985,7415,8961,9865,10066,11201,11777,12745,15265,15625,
294,348,626,815,1226,2381,3726,4106,6505,6986,7416,8962,9866,10067,11202,11778,12746,15266,15626,
295,349,627,816,1227,2382,3727,4107,6506,6987,7417,8963,9867,10068,11203,11779,12747,15267,15627,
296,350,628,817,1228,2383,3728,4108,6507,6988,7418,8964,9868,10069,11204,11780,12748,15268,15628,
297,351,629,818,1229,2384,3729,4109,6508,6989,7419,8965,9869,10070,11205,11781,12749,15269,15629,
298,352,630,819,1230,2385,3730,4110,6509,6990,7420,8966,9870,10071,11206,11782,12750,15270,15630,
299,353,631,820,1231,2386,3731,4111,6510,6991,7421,8967,9871,10072,11207,11783,12751,15271,15631,
300,354,632,821,1232,2387,3732,4112,6511,6992,7422,8968,9872,10073,11208,11784,12752,15272,15632,
301,355,633,822,1233,2388,3733,4113,6512,6993,7423,8969,9873,10074,11209,11785,12753,15273,15633,
302,356,634,823,1234,2389,3734,4114,6513,6994,7424,8970,9874,10075,11210,11786,12754,15274,15634,
303,357,635,824,1235,2390,3735,4115,6514,6995,7425,8971,9875,10076,11211,11787,12755,15275,15635,
304,358,636,825,1236,2391,3736,4116,6515,6996,7426,8972,9876,10077,11212,11788,12756,15276,15636,
305,359,637,826,1237,2392,3737,4117,6516,6997,7427,8973,9877,10078,11213,11789,12757,15277,15637,
0,306,638,827,1238,2393,3738,4118,6517,6998,7428,8974,9878,10079,11214,11790,12758,15278,15638,
1,307,639,828,1239,2394,3739,4119,6518,6999,7429,8975,9720,9879,11215,11791,12759,15279,15639,
2,308,640,829,1240,2395,3740,4120,6519,7000,7430,8976,9721,9880,11216,11792,12760,15280,15640,
3,309,641,830,1241,2396,3741,4121,6520,7001,7431,8977,9722,9881,11217,11793,12761,15281,15641,
4,310,642,831,1242,2397,3742,4122,6521,7002,7432,8978,9723,9882,11218,11794,12762,15282,15642,
5,311,643,832,1243,2398,3743,4123,6522,7003,7433,8979,9724,9883,11219,11795,12763,15283,15643,
6,312,644,833,1244,2399,3744,4124,6523,7004,7434,8980,9725,9884,11220,11796,12764,15284,15644,
7,313,645,834,1245,2400,3745,4125,6524,7005,7435,8981,9726,9885,11221,11797,12765,15285,15645,
8,314,646,835,1246,2401,3746,4126,6525,7006,7436,8982,9727,9886,11222,11798,12766,15286,15646,
9,315,647,836,1247,2402,3747,4127,6526,7007,7437,8983,9728,9887,11223,11799,12767,15287,15647,
10,316,648,837,1248,2403,3748,4128,6527,7008,7438,8984,9729,9888,11224,11800,12768,15288,15648,
11,317,649,838,1249,2404,3749,4129,6528,7009,7439,8985,9730,9889,11225,11801,12769,15289,15649,
12,318,650,839,1250,2405,3750,4130,6529,7010,7440,8986,9731,9890,11226,11802,12770,15290,15650,
13,319,651,840,1251,2406,3751,4131,6530,7011,7441,8987,9732,9891,11227,11803,12771,15291,15651,
14,320,652,841,1252,2407,3752,4132,6531,7012,7442,8988,9733,9892,11228,11804,12772,15292,15652,
15,321,653,842,1253,2408,3753,4133,6532,7013,7443,8989,9734,9893,11229,11805,12773,15293,15653,
16,322,654,843,1254,2409,3754,4134,6533,7014,7444,8990,9735,9894,11230,11806,12774,15294,15654,
17,323,655,844,1255,2410,3755,4135,6534,7015,7445,8991,9736,9895,11231,11807,12775,15295,15655,
18,324,656,845,1256,2411,3756,4136,6535,7016,7446,8992,9737,9896,11232,11808,12776,15296,15656,
19,325,657,846,1257,2412,3757,4137,6536,7017,7447,8993,9738,9897,11233,11809,12777,15297,15657,
20,326,658,847,1258,2413,3758,4138,6537,7018,7448,8994,9739,9898,11234,11810,12778,15298,15658,
21,327,659,848,1259,2414,3759,4139,6538,7019,7449,8995,9740,9899,11235,11811,12779,15299,15659,
22,328,660,849,1260,2415,3760,4140,6539,7020,7450,8996,9741,9900,11236,11812,12780,15300,15660,
23,329,661,850,1261,2416,3761,4141,6540,7021,7451,8997,9742,9901,11237,11813,12781,15301,15661,
24,330,662,851,1262,2417,3762,4142,6541,7022,7452,8998,9743,9902,11238,11814,12782,15302,15662,
25,331,663,852,1263,2418,3763,4143,6542,7023,7453,8999,9744,9903,11239,11815,12783,15303,15663,
26,332,664,853,1264,2419,3764,4144,6543,7024,7454,8640,9745,9904,11240,11816,12784,15304,15664,
27,333,665,854,1265,2420,3765,4145,6544,7025,7455,8641,9746,9905,11241,11817,12785,15305,15665,
28,334,666,855,1266,2421,3766,4146,6545,7026,7456,8642,9747,9906,11242,11818,12786,15306,15666,
29,335,667,856,1267,2422,3767,4147,6546,7027,7457,8643,9748,9907,11243,11819,12787,15307,15667,
30,336,668,857,1268,2423,3768,4148,6547,7028,7458,8644,9749,9908,11244,11820,12788,15308,15668,
31,337,669,858,1269,2424,3769,4149,6548,7029,7459,8645,9750,9909,11245,11821,12789,15309,15669,
32,338,670,859,1270,2425,3770,4150,6549,7030,7460,8646,9751,9910,11246,11822,12790,15310,15670,
33,339,671,860,1271,2426,3771,4151,6550,7031,7461,8647,9752,9911,11247,11823,12791,15311,15671,
34,340,672,861,1272,2427,3772,4152,6551,7032,7462,8648,9753,9912,11248,11824,12792,15312,15672,
35,341,673,862,1273,2428,3773,4153,6552,7033,7463,8649,9754,9913,11249,11825,12793,15313,15673,
36,342,674,863,1274,2429,3774,4154,6553,7034,7464,8650,9755,9914,11250,11826,12794,15314,15674,
37,343,675,864,1275,2430,3775,4155,6554,7035,7465,8651,9756,9915,11251,11827,12795,15315,15675,
38,344,676,865,1276,2431,3776,4156,6555,7036,7466,8652,9757,9916,11252,11828,12796,15316,15676,
39,345,677,866,1277,2432,3777,4157,6556,7037,7467,8653,9758,9917,11253,11829,12797,15317,15677,
40,346,678,867,1278,2433,3778,4158,6557,7038,7468,8654,9759,9918,11254,11830,12798,15318,15678,
41,347,679,868,1279,2434,3779,4159,6558,7039,7469,8655,9760,9919,11255,11831,12799,15319,15679,
42,348,680,869,1280,2435,3780,4160,6559,7040,7470,8656,9761,9920,11256,11832,12800,15320,15680,
43,349,681,870,1281,2436,3781,4161,6560,7041,7471,8657,9762,9921,11257,11833,12801,15321,15681,
44,350,682,871,1282,2437,3782,4162,6561,7042,7472,8658,9763,9922,11258,11834,12802,15322,15682,
45,351,683,872,1283,2438,3783,4163,6562,7043,7473,8659,9764,9923,11259,11835,12803,15323,15683,
46,352,684,873,1284,2439,3784,4164,6563,7044,7474,8660,9765,9924,11260,11836,12804,15324,15684,
47,353,685,874,1285,2440,3785,4165,6564,7045,7475,8661,9766,9925,11261,11837,12805,15325,15685,
48,354,686,875,1286,2441,3786,4166,6565,7046,7476,8662,9767,9926,11262,11838,12806,15326,15686,
49,355,687,876,1287,2442,3787,4167,6566,7047,7477,8663,9768,9927,11263,11839,12807,15327,15687,
50,356,688,877,1288,2443,3788,4168,6567,7048,7478,8664,9769,9928,11264,11840,12808,15328,15688,
51,357,689,878,1289,2444,3789,4169,6568,7049,7479,8665,9770,9929,11265,11841,12809,15329,15689,
52,358,690,879,1290,2445,3790,4170,6569,7050,7480,8666,9771,9930,11266,11842,12810,15330,15690,
53,359,691,880,1291,2446,3791,4171,6570,7051,7481,8667,9772,9931,11267,11843,12811,15331,15691,
0,54,692,881,1292,2447,3792,4172,6571,7052,7482,8668,9773,9932,11268,11844,12812,15332,15692,
1,55,693,882,1293,2448,3793,4173,6572,7053,7483,8669,9774,9933,11269,11845,12813,15333,15693,
2,56,694,883,1294,2449,3794,4174,6573,7054,7484,8670,9775,9934,11270,11846,12814,15334,15694,
3,57,695,884,1295,2450,3795,4175,6574,7055,7485,8671,9776,9935,11271,11847,12815,15335,15695,
4,58,696,885,1296,2451,3796,4176,6575,7056,7486,8672,9777,9936,11272,11848,12816,15336,15696,
5,59,697,886,1297,2452,3797,4177,6576,7057,7487,8673,9778,9937,11273,11849,12817,15337,15697,
6,60,698,887,1298,2453,3798,4178,6577,7058,7488,8674,9779,9938,11274,11850,12818,15338,15698,
7,61,699,888,1299,2454,3799,4179,6578,7059,7489,8675,9780,9939,11275,11851,12819,15339,15699,
8,62,700,889,1300,2455,3800,4180,6579,7060,7490,8676,9781,9940,11276,11852,12820,15340,15700,
9,63,701,890,1301,2456,3801,4181,6580,7061,7491,8677,9782,9941,11277,11853,12821,15341,15701,
10,64,702,891,1302,2457,3802,4182,6581,7062,7492,8678,9783,9942,11278,11854,12822,15342,15702,
11,65,703,892,1303,2458,3803,4183,6582,7063,7493,8679,9784,9943,11279,11855,12823,15343,15703,
12,66,704,893,1304,2459,3804,4184,6583,7064,7494,8680,9785,9944,11280,11856,12824,15344,15704,
13,67,705,894,1305,2460,3805,4185,6584,7065,7495,8681,9786,9945,11281,11857,12825,15345,15705,
14,68,706,895,1306,2461,3806,4186,6585,7066,7496,8682,9787,9946,11282,11858,12826,15346,15706,
15,69,707,896,1307,2462,3807,4187,6586,7067,7497,8683,9788,9947,11283,11859,12827,15347,15707,
16,70,708,897,1308,2463,3808,4188,6587,7068,7498,8684,9789,9948,11284,11860,12828,15348,15708,
17,71,709,898,1309,2464,3809,4189,6588,7069,7499,8685,9790,9949,11285,11861,12829,15349,15709,
18,72,710,899,1310,2465,3810,4190,6589,7070,7500,8686,9791,9950,11286,11862,12830,15350,15710,
19,73,711,900,1311,2466,3811,4191,6590,7071,7501,8687,9792,9951,11287,11863,12831,15351,15711,
20,74,712,901,1312,2467,3812,4192,6591,7072,7502,8688,9793,9952,11288,11864,12832,15352,15712,
21,75,713,902,1313,2468,3813,4193,6592,7073,7503,8689,9794,9953,11289,11865,12833,15353,15713,
22,76,714,903,1314,2469,3814,4194,6593,7074,7504,8690,9795,9954,11290,11866,12834,15354,15714,
23,77,715,904,1315,2470,3815,4195,6594,7075,7505,8691,9796,9955,11291,11867,12835,15355,15715,
24,78,716,905,1316,2471,3816,4196,6595,7076,7506,8692,9797,9956,11292,11868,12836,15356,15716,
25,79,717,906,1317,2472,3817,4197,6596,7077,7507,8693,9798,9957,11293,11869,12837,15357,15717,
26,80,718,907,1318,2473,3818,4198,6597,7078,7508,8694,9799,9958,11294,11870,12838,15358,15718,
27,81,719,908,1319,2474,3819,4199,6598,7079,7509,8695,9800,9959,11295,11871,12839,15359,15719,
28,82,360,909,1320,2475,3820,4200,6599,7080,7510,8696,9801,9960,11296,11872,12840,15360,15720,
29,83,361,910,1321,2476,3821,4201,6600,7081,7511,8697,9802,9961,11297,11873,12841,15361,15721,
30,84,362,911,1322,2477,3822,4202,6601,7082,7512,8698,9803,9962,11298,11874,12842,15362,15722,
31,85,363,912,1323,2478,3823,4203,6602,7083,7513,8699,9804,9963,11299,11875,12843,15363,15723,
32,86,364,913,1324,2479,3824,4204,6603,7084,7514,8700,9805,9964,11300,11876,12844,15364,15724,
33,87,365,914,1325,2480,3825,4205,6604,7085,7515,8701,9806,9965,11301,11877,12845,15365,15725,
34,88,366,915,1326,2481,3826,4206,6605,7086,7516,8702,9807,9966,11302,11878,12846,15366,15726,
35,89,367,916,1327,2482,3827,4207,6606,7087,7517,8703,9808,9967,11303,11879,12847,15367,15727,
36,90,368,917,1328,2483,3828,4208,6607,7088,7518,8704,9809,9968,11304,11520,12848,15368,15728,
37,91,369,918,1329,2484,3829,4209,6608,7089,7519,8705,9810,9969,11305,11521,12849,15369,15729,
38,92,370,919,1330,2485,3830,4210,6609,7090,7520,8706,9811,9970,11306,11522,12850,15370,15730,
39,93,371,920,1331,2486,3831,4211,6610,7091,7521,8707,9812,9971,11307,11523,12851,15371,15731,
40,94,372,921,1332,2487,3832,4212,6611,7092,7522,8708,9813,9972,11308,11524,12852,15372,15732,
41,95,373,922,1333,2488,3833,4213,6612,7093,7523,8709,9814,9973,11309,11525,12853,15373,15733,
42,96,374,923,1334,2489,3834,4214,6613,7094,7524,8710,9815,9974,11310,11526,12854,15374,15734,
43,97,375,924,1335,2490,3835,4215,6614,7095,7525,8711,9816,9975,11311,11527,12855,15375,15735,
44,98,376,925,1336,2491,3836,4216,6615,7096,7526,8712,9817,9976,11312,11528,12856,15376,15736,
45,99,377,926,1337,2492,3837,4217,6616,7097,7527,8713,9818,9977,11313,11529,12857,15377,15737,
46,100,378,927,1338,2493,3838,4218,6617,7098,7528,8714,9819,9978,11314,11530,12858,15378,15738,
47,101,379,928,1339,2494,3839,4219,6618,7099,7529,8715,9820,9979,11315,11531,12859,15379,15739,
48,102,380,929,1340,2495,3840,4220,6619,7100,7530,8716,9821,9980,11316,11532,12860,15380,15740,
49,103,381,930,1341,2496,3841,4221,6620,7101,7531,8717,9822,9981,11317,11533,12861,15381,15741,
50,104,382,931,1342,2497,3842,4222,6621,7102,7532,8718,9823,9982,11318,11534,12862,15382,15742,
51,105,383,932,1343,2498,3843,4223,6622,7103,7533,8719,9824,9983,11319,11535,12863,15383,15743,
52,106,384,933,1344,2499,3844,4224,6623,7104,7534,8720,9825,9984,11320,11536,12864,15384,15744,
53,107,385,934,1345,2500,3845,4225,6624,7105,7535,8721,9826,9985,11321,11537,12865,15385,15745,
54,108,386,935,1346,2501,3846,4226,6625,7106,7536,8722,9827,9986,11322,11538,12866,15386,15746,
55,109,387,936,1347,2502,3847,4227,6626,7107,7537,8723,9828,9987,11323,11539,12867,15387,15747,
56,110,388,937,1348,2503,3848,4228,6627,7108,7538,8724,9829,9988,11324,11540,12868,15388,15748,
57,111,389,938,1349,2504,3849,4229,6628,7109,7539,8725,9830,9989,11325,11541,12869,15389,15749,
58,112,390,939,1350,2505,3850,4230,6629,7110,7540,8726,9831,9990,11326,11542,12870,15390,15750,
59,113,391,940,1351,2506,3851,4231,6630,7111,7541,8727,9832,9991,11327,11543,12871,15391,15751,
60,114,392,941,1352,2507,3852,4232,6631,7112,7542,8728,9833,9992,11328,11544,12872,15392,15752,
61,115,393,942,1353,2508,3853,4233,6632,7113,7543,8729,9834,9993,11329,11545,12873,15393,15753,
62,116,394,943,1354,2509,3854,4234,6633,7114,7544,8730,9835,9994,11330,11546,12874,15394,15754,
63,117,395,944,1355,2510,3855,4235,6634,7115,7545,8731,9836,9995,11331,11547,12875,15395,15755,
64,118,396,945,1356,2511,3856,4236,6635,7116,7546,8732,9837,9996,11332,11548,12876,15396,15756,
65,119,397,946,1357,2512,3857,4237,6636,7117,7547,8733,9838,9997,11333,11549,12877,15397,15757,
66,120,398,947,1358,2513,3858,4238,6637,7118,7548,8734,9839,9998,11334,11550,12878,15398,15758,
67,121,399,948,1359,2514,3859,4239,6638,7119,7549,8735,9840,9999,11335,11551,12879,15399,15759,
68,122,400,949,1360,2515,3860,4240,6639,7120,7550,8736,9841,10000,11336,11552,12880,15400,15760,
69,123,401,950,1361,2516,3861,4241,6640,7121,7551,8737,9842,10001,11337,11553,12881,15401,15761,
70,124,402,951,1362,2517,3862,4242,6641,7122,7552,8738,9843,10002,11338,11554,12882,15402,15762,
71,125,403,952,1363,2518,3863,4243,6642,7123,7553,8739,9844,10003,11339,11555,12883,15403,15763,
72,126,404,953,1364,2519,3864,4244,6643,7124,7554,8740,9845,10004,11340,11556,12884,15404,15764,
73,127,405,954,1365,2160,3865,4245,6644,7125,7555,8741,9846,10005,11341,11557,12885,15405,15765,
74,128,406,955,1366,2161,3866,4246,6645,7126,7556,8742,9847,10006,11342,11558,12886,15406,15766,
75,129,407,956,1367,2162,3867,4247,6646,7127,7557,8743,9848,10007,11343,11559,12887,15407,15767,
76,130,408,957,1368,2163,3868,4248,6647,7128,7558,8744,9849,10008,11344,11560,12888,15408,15768,
77,131,409,958,1369,2164,3869,4249,6648,7129,7559,8745,9850,10009,11345,11561,12889,15409,15769,
78,132,410,959,1370,2165,3870,4250,6649,7130,7200,8746,9851,10010,11346,11562,12890,15410,15770,
79,133,411,960,1371,2166,3871,4251,6650,7131,7201,8747,9852,10011,11347,11563,12891,15411,15771,
80,134,412,961,1372,2167,3872,4252,6651,7132,7202,8748,9853,10012,11348,11564,12892,15412,15772,
81,135,413,962,1373,2168,3873,4253,6652,7133,7203,8749,9854,10013,11349,11565,12893,15413,15773,
82,136,414,963,1374,2169,3874,4254,6653,7134,7204,8750,9855,10014,11350,11566,12894,15414,15774,
83,137,415,964,1375,2170,3875,4255,6654,7135,7205,8751,9856,10015,11351,11567,12895,15415,15775,
84,138,416,965,1376,2171,3876,4256,6655,7136,7206,8752,9857,10016,11352,11568,12896,15416,15776,
85,139,417,966,1377,2172,3877,4257,6656,7137,7207,8753,9858,10017,11353,11569,12897,15417,15777,
86,140,418,967,1378,2173,3878,4258,6657,7138,7208,8754,9859,10018,11354,11570,12898,15418,15778,
87,141,419,968,1379,2174,3879,4259,6658,7139,7209,8755,9860,10019,11355,11571,12899,15419,15779,
88,142,420,969,1380,2175,3880,4260,6659,7140,7210,8756,9861,10020,11356,11572,12900,15420,15780,
89,143,421,970,1381,2176,3881,4261,6660,7141,7211,8757,9862,10021,11357,11573,12901,15421,15781,
90,144,422,971,1382,2177,3882,4262,6661,7142,7212,8758,9863,10022,11358,11574,12902,15422,15782,
91,145,423,972,1383,2178,3883,4263,6662,7143,7213,8759,9864,10023,11359,11575,12903,15423,15783,
92,146,424,973,1384,2179,3884,4264,6663,7144,7214,8760,9865,10024,11360,11576,12904,15424,15784,
93,147,425,974,1385,2180,3885,4265,6664,7145,7215,8761,9866,10025,11361,11577,12905,15425,15785,
94,148,426,975,1386,2181,3886,4266,6665,7146,7216,8762,9867,10026,11362,11578,12906,15426,15786,
95,149,427,976,1387,2182,3887,4267,6666,7147,7217,8763,9868,10027,11363,11579,12907,15427,15787,
96,150,428,977,1388,2183,3888,4268,6667,7148,7218,8764,9869,10028,11364,11580,12908,15428,15788,
97,151,429,978,1389,2184,3889,4269,6668,7149,7219,8765,9870,10029,11365,11581,12909,15429,15789,
98,152,430,979,1390,2185,3890,4270,6669,7150,7220,8766,9871,10030,11366,11582,12910,15430,15790,
99,153,431,980,1391,2186,3891,4271,6670,7151,7221,8767,9872,10031,11367,11583,12911,15431,15791,
100,154,432,981,1392,2187,3892,4272,6671,7152,7222,8768,9873,10032,11368,11584,12912,15432,15792,
101,155,433,982,1393,2188,3893,4273,6672,7153,7223,8769,9874,10033,11369,11585,12913,15433,15793,
102,156,434,983,1394,2189,3894,4274,6673,7154,7224,8770,9875,10034,11370,11586,12914,15434,15794,
103,157,435,984,1395,2190,3895,4275,6674,7155,7225,8771,9876,10035,11371,11587,12915,15435,15795,
104,158,436,985,1396,2191,3896,4276,6675,7156,7226,8772,9877,10036,11372,11588,12916,15436,15796,
105,159,437,986,1397,2192,3897,4277,6676,7157,7227,8773,9878,10037,11373,11589,12917,15437,15797,
106,160,438,987,1398,2193,3898,4278,6677,7158,7228,8774,9879,10038,11374,11590,12918,15438,15798,
107,161,439,988,1399,2194,3899,4279,6678,7159,7229,8775,9880,10039,11375,11591,12919,15439,15799,
108,162,440,989,1400,2195,3900,4280,6679,7160,7230,8776,9881,10040,11376,11592,12920,15440,15800,
109,163,441,990,1401,2196,3901,4281,6680,7161,7231,8777,9882,10041,11377,11593,12921,15441,15801,
110,164,442,991,1402,2197,3902,4282,6681,7162,7232,8778,9883,10042,11378,11594,12922,15442,15802,
111,165,443,992,1403,2198,3903,4283,6682,7163,7233,8779,9884,10043,11379,11595,12923,15443,15803,
112,166,444,993,1404,2199,3904,4284,6683,7164,7234,8780,9885,10044,11380,11596,12924,15444,15804,
113,167,445,994,1405,2200,3905,4285,6684,7165,7235,8781,9886,10045,11381,11597,12925,15445,15805,
114,168,446,995,1406,2201,3906,4286,6685,7166,7236,8782,9887,10046,11382,11598,12926,15446,15806,
115,169,447,996,1407,2202,3907,4287,6686,7167,7237,8783,9888,10047,11383,11599,12927,15447,15807,
116,170,448,997,1408,2203,3908,4288,6687,7168,7238,8784,9889,10048,11384,11600,12928,15448,15808,
117,171,449,998,1409,2204,3909,4289,6688,7169,7239,8785,9890,10049,11385,11601,12929,15449,15809,
118,172,450,999,1410,2205,3910,4290,6689,7170,7240,8786,9891,10050,11386,11602,12930,15450,15810,
119,173,451,1000,1411,2206,3911,4291,6690,7171,7241,8787,9892,10051,11387,11603,12931,15451,15811,
120,174,452,1001,1412,2207,3912,4292,6691,7172,7242,8788,9893,10052,11388,11604,12932,15452,15812,
121,175,453,1002,1413,2208,3913,4293,6692,7173,7243,8789,9894,10053,11389,11605,12933,15453,15813,
122,176,454,1003,1414,2209,3914,4294,6693,7174,7244,8790,9895,10054,11390,11606,12934,15454,15814,
123,177,455,1004,1415,2210,3915,4295,6694,7175,7245,8791,9896,10055,11391,11607,12935,15455,15815,
124,178,456,1005,1416,2211,3916,4296,6695,7176,7246,8792,9897,10056,11392,11608,12936,15456,15816,
125,179,457,1006,1417,2212,3917,4297,6696,7177,7247,8793,9898,10057,11393,11609,12937,15457,15817,
126,180,458,1007,1418,2213,3918,4298,6697,7178,7248,8794,9899,10058,11394,11610,12938,15458,15818,
127,181,459,1008,1419,2214,3919,4299,6698,7179,7249,8795,9900,10059,11395,11611,12939,15459,15819,
128,182,460,1009,1420,2215,3920,4300,6699,7180,7250,8796,9901,10060,11396,11612,12940,15460,15820,
129,183,461,1010,1421,2216,3921,4301,6700,7181,7251,8797,9902,10061,11397,11613,12941,15461,15821,
130,184,462,1011,1422,2217,3922,4302,6701,7182,7252,8798,9903,10062,11398,11614,12942,15462,15822,
131,185,463,1012,1423,2218,3923,4303,6702,7183,7253,8799,9904,10063,11399,11615,12943,15463,15823,
132,186,464,1013,1424,2219,3924,4304,6703,7184,7254,8800,9905,10064,11400,11616,12944,15464,15824,
133,187,465,1014,1425,2220,3925,4305,6704,7185,7255,8801,9906,10065,11401,11617,12945,15465,15825,
134,188,466,1015,1426,2221,3926,4306,6705,7186,7256,8802,9907,10066,11402,11618,12946,15466,15826,
135,189,467,1016,1427,2222,3927,4307,6706,7187,7257,8803,9908,10067,11403,11619,12947,15467,15827,
136,190,468,1017,1428,2223,3928,4308,6707,7188,7258,8804,9909,10068,11404,11620,12948,15468,15828,
137,191,469,1018,1429,2224,3929,4309,6708,7189,7259,8805,9910,10069,11405,11621,12949,15469,15829,
138,192,470,1019,1430,2225,3930,4310,6709,7190,7260,8806,9911,10070,11406,11622,12950,15470,15830,
139,193,471,1020,1431,2226,3931,4311,6710,7191,7261,8807,9912,10071,11407,11623,12951,15471,15831,
140,194,472,1021,1432,2227,3932,4312,6711,7192,7262,8808,9913,10072,11408,11624,12952,15472,15832,
141,195,473,1022,1433,2228,3933,4313,6712,7193,7263,8809,9914,10073,11409,11625,12953,15473,15833,
142,196,474,1023,1434,2229,3934,4314,6713,7194,7264,8810,9915,10074,11410,11626,12954,15474,15834,
143,197,475,1024,1435,2230,3935,4315,6714,7195,7265,8811,9916,10075,11411,11627,12955,15475,15835,
144,198,476,1025,1436,2231,3936,4316,6715,7196,7266,8812,9917,10076,11412,11628,12956,15476,15836,
145,199,477,1026,1437,2232,3937,4317,6716,7197,7267,8813,9918,10077,11413,11629,12957,15477,15837,
146,200,478,1027,1438,2233,3938,4318,6717,7198,7268,8814,9919,10078,11414,11630,12958,15478,15838,
147,201,479,1028,1439,2234,3939,4319,6718,7199,7269,8815,9920,10079,11415,11631,12959,15479,15839,
291,415,1440,1863,3223,4320,5304,5767,7200,9047,10080,10378,11727,12482,12960,15480,15840,
292,416,1441,1864,3224,4321,5305,5768,7201,9048,10081,10379,11728,12483,12961,15481,15841,
293,417,1442,1865,3225,4322,5306,5769,7202,9049,10082,10380,11729,12484,12962,15482,15842,
294,418,1443,1866,3226,4323,5307,5770,7203,9050,10083,10381,11730,12485,12963,15483,15843,
295,419,1444,1867,3227,4324,5308,5771,7204,9051,10084,10382,11731,12486,12964,15484,15844,
296,420,1445,1868,3228,4325,5309,5772,7205,9052,10085,10383,11732,12487,12965,15485,15845,
297,421,1446,1869,3229,4326,5310,5773,7206,9053,10086,10384,11733,12488,12966,15486,15846,
298,422,1447,1870,3230,4327,5311,5774,7207,9054,10087,10385,11734,12489,12967,15487,15847,
299,423,1448,1871,3231,4328,5312,5775,7208,9055,10088,10386,11735,12490,12968,15488,15848,
300,424,1449,1872,3232,4329,5313,5776,7209,9056,10089,10387,11736,12491,12969,15489,15849,
301,425,1450,1873,3233,4330,5314,5777,7210,9057,10090,10388,11737,12492,12970,15490,15850,
302,426,1451,1874,3234,4331,5315,5778,7211,9058,10091,10389,11738,12493,12971,15491,15851,
303,427,1452,1875,3235,4332,5316,5779,7212,9059,10092,10390,11739,12494,12972,15492,15852,
304,428,1453,1876,3236,4333,5317,5780,7213,9060,10093,10391,11740,12495,12973,15493,15853,
305,429,1454,1877,3237,4334,5318,5781,7214,9061,10094,10392,11741,12496,12974,15494,15854,
306,430,1455,1878,3238,4335,5319,5782,7215,9062,10095,10393,11742,12497,12975,15495,15855,
307,431,1456,1879,3239,4336,5320,5783,7216,9063,10096,10394,11743,12498,12976,15496,15856,
308,432,1457,1880,2880,4337,5321,5784,7217,9064,10097,10395,11744,12499,12977,15497,15857,
309,433,1458,1881,2881,4338,5322,5785,7218,9065,10098,10396,11745,12500,12978,15498,15858,
310,434,1459,1882,2882,4339,5323,5786,7219,9066,10099,10397,11746,12501,12979,15499,15859,
311,435,1460,1883,2883,4340,5324,5787,7220,9067,10100,10398,11747,12502,12980,15500,15860,
312,436,1461,1884,2884,4341,5325,5788,7221,9068,10101,10399,11748,12503,12981,15501,15861,
313,437,1462,1885,2885,4342,5326,5789,7222,9069,10102,10400,11749,12504,12982,15502,15862,
314,438,1463,1886,2886,4343,5327,5790,7223,9070,10103,10401,11750,12505,12983,15503,15863,
315,439,1464,1887,2887,4344,5328,5791,7224,9071,10104,10402,11751,12506,12984,15504,15864,
316,440,1465,1888,2888,4345,5329,5792,7225,9072,10105,10403,11752,12507,12985,15505,15865,
317,441,1466,1889,2889,4346,5330,5793,7226,9073,10106,10404,11753,12508,12986,15506,15866,
318,442,1467,1890,2890,4347,5331,5794,7227,9074,10107,10405,11754,12509,12987,15507,15867,
319,443,1468,1891,2891,4348,5332,5795,7228,9075,10108,10406,11755,12510,12988,15508,15868,
320,444,1469,1892,2892,4349,5333,5796,7229,9076,10109,10407,11756,12511,12989,15509,15869,
321,445,1470,1893,2893,4350,5334,5797,7230,9077,10110,10408,11757,12512,12990,15510,15870,
322,446,1471,1894,2894,4351,5335,5798,7231,9078,10111,10409,11758,12513,12991,15511,15871,
323,447,1472,1895,2895,4352,5336,5799,7232,9079,10112,10410,11759,12514,12992,15512,15872,
324,448,1473,1896,2896,4353,5337,5800,7233,9080,10113,10411,11760,12515,12993,15513,15873,
325,449,1474,1897,2897,4354,5338,5801,7234,9081,10114,10412,11761,12516,12994,15514,15874,
326,450,1475,1898,2898,4355,5339,5802,7235,9082,10115,10413,11762,12517,12995,15515,15875,
327,451,1476,1899,2899,4356,5340,5803,7236,9083,10116,10414,11763,12518,12996,15516,15876,
328,452,1477,1900,2900,4357,5341,5804,7237,9084,10117,10415,11764,12519,12997,15517,15877,
329,453,1478,1901,2901,4358,5342,5805,7238,9085,10118,10416,11765,12520,12998,15518,15878,
330,454,1479,1902,2902,4359,5343,5806,7239,9086,10119,10417,11766,12521,12999,15519,15879,
331,455,1480,1903,2903,4360,5344,5807,7240,9087,10120,10418,11767,12522,13000,15520,15880,
332,456,1481,1904,2904,4361,5345,5808,7241,9088,10121,10419,11768,12523,13001,15521,15881,
333,457,1482,1905,2905,4362,5346,5809,7242,9089,10122,10420,11769,12524,13002,15522,15882,
334,458,1483,1906,2906,4363,5347,5810,7243,9090,10123,10421,11770,12525,13003,15523,15883,
335,459,1484,1907,2907,4364,5348,5811,7244,9091,10124,10422,11771,12526,13004,15524,15884,
336,460,1485,1908,2908,4365,5349,5812,7245,9092,10125,10423,11772,12527,13005,15525,15885,
337,461,1486,1909,2909,4366,5350,5813,7246,9093,10126,10424,11773,12528,13006,15526,15886,
338,462,1487,1910,2910,4367,5351,5814,7247,9094,10127,10425,11774,12529,13007,15527,15887,
339,463,1488,1911,2911,4368,5352,5815,7248,9095,10128,10426,11775,12530,13008,15528,15888,
340,464,1489,1912,2912,4369,5353,5816,7249,9096,10129,10427,11776,12531,13009,15529,15889,
341,465,1490,1913,2913,4370,5354,5817,7250,9097,10130,10428,11777,12532,13010,15530,15890,
342,466,1491,1914,2914,4371,5355,5818,7251,9098,10131,10429,11778,12533,13011,15531,15891,
343,467,1492,1915,2915,4372,5356,5819,7252,9099,10132,10430,11779,12534,13012,15532,15892,
344,468,1493,1916,2916,4373,5357,5820,7253,9100,10133,10431,11780,12535,13013,15533,15893,
345,469,1494,1917,2917,4374,5358,5821,7254,9101,10134,10432,11781,12536,13014,15534,15894,
346,470,1495,1918,2918,4375,5359,5822,7255,9102,10135,10433,11782,12537,13015,15535,15895,
347,471,1496,1919,2919,4376,5360,5823,7256,9103,10136,10434,11783,12538,13016,15536,15896,
348,472,1497,1920,2920,4377,5361,5824,7257,9104,10137,10435,11784,12539,13017,15537,15897,
349,473,1498,1921,2921,4378,5362,5825,7258,9105,10138,10436,11785,12540,13018,15538,15898,
350,474,1499,1922,2922,4379,5363,5826,7259,9106,10139,10437,11786,12541,13019,15539,15899,
351,475,1500,1923,2923,4380,5364,5827,7260,9107,10140,10438,11787,12542,13020,15540,15900,
352,476,1501,1924,2924,4381,5365,5828,7261,9108,10141,10439,11788,12543,13021,15541,15901,
353,477,1502,1925,2925,4382,5366,5829,7262,9109,10080,10142,11789,12544,13022,15542,15902,
354,478,1503,1926,2926,4383,5367,5830,7263,9110,10081,10143,11790,12545,13023,15543,15903,
355,479,1504,1927,2927,4384,5368,5831,7264,9111,10082,10144,11791,12546,13024,15544,15904,
356,480,1505,1928,2928,4385,5369,5832,7265,9112,10083,10145,11792,12547,13025,15545,15905,
357,481,1506,1929,2929,4386,5370,5833,7266,9113,10084,10146,11793,12548,13026,15546,15906,
358,482,1507,1930,2930,4387,5371,5834,7267,9114,10085,10147,11794,12549,13027,15547,15907,
359,483,1508,1931,2931,4388,5372,5835,7268,9115,10086,10148,11795,12550,13028,15548,15908,
0,484,1509,1932,2932,4389,5373,5836,7269,9116,10087,10149,11796,12551,13029,15549,15909,
1,485,1510,1933,2933,4390,5374,5837,7270,9117,10088,10150,11797,12552,13030,15550,15910,
2,486,1511,1934,2934,4391,5375,5838,7271,9118,10089,10151,11798,12553,13031,15551,15911,
3,487,1512,1935,2935,4392,5376,5839,7272,9119,10090,10152,11799,12554,13032,15552,15912,
4,488,1513,1936,2936,4393,5377,5840,7273,9120,10091,10153,11800,12555,13033,15553,15913,
5,489,1514,1937,2937,4394,5378,5841,7274,9121,10092,10154,11801,12556,13034,15554,15914,
6,490,1515,1938,2938,4395,5379,5842,7275,9122,10093,10155,11802,12557,13035,15555,15915,
7,491,1516,1939,2939,4396,5380,5843,7276,9123,10094,10156,11803,12558,13036,15556,15916,
8,492,1517,1940,2940,4397,5381,5844,7277,9124,10095,10157,11804,12559,13037,15557,15917,
9,493,1518,1941,2941,4398,5382,5845,7278,9125,10096,10158,11805,12560,13038,15558,15918,
10,494,1519,1942,2942,4399,5383,5846,7279,9126,10097,10159,11806,12561,13039,15559,15919,
11,495,1520,1943,2943,4400,5384,5847,7280,9127,10098,10160,11807,12562,13040,15560,15920,
12,496,1521,1944,2944,4401,5385,5848,7281,9128,10099,10161,11808,12563,13041,15561,15921,
13,497,1522,1945,2945,4402,5386,5849,7282,9129,10100,10162,11809,12564,13042,15562,15922,
14,498,1523,1946,2946,4403,5387,5850,7283,9130,10101,10163,11810,12565,13043,15563,15923,
15,499,1524,1947,2947,4404,5388,5851,7284,9131,10102,10164,11811,12566,13044,15564,15924,
16,500,1525,1948,2948,4405,5389,5852,7285,9132,10103,10165,11812,12567,13045,15565,15925,
17,501,1526,1949,2949,4406,5390,5853,7286,9133,10104,10166,11813,12568,13046,15566,15926,
18,502,1527,1950,2950,4407,5391,5854,7287,9134,10105,10167,11814,12569,13047,15567,15927,
19,503,1528,1951,2951,4408,5392,5855,7288,9135,10106,10168,11815,12570,13048,15568,15928,
20,504,1529,1952,2952,4409,5393,5856,7289,9136,10107,10169,11816,12571,13049,15569,15929,
21,505,1530,1953,2953,4410,5394,5857,7290,9137,10108,10170,11817,12572,13050,15570,15930,
22,506,1531,1954,2954,4411,5395,5858,7291,9138,10109,10171,11818,12573,13051,15571,15931,
23,507,1532,1955,2955,4412,5396,5859,7292,9139,10110,10172,11819,12574,13052,15572,15932,
24,508,1533,1956,2956,4413,5397,5860,7293,9140,10111,10173,11820,12575,13053,15573,15933,
25,509,1534,1957,2957,4414,5398,5861,7294,9141,10112,10174,11821,12576,13054,15574,15934,
26,510,1535,1958,2958,4415,5399,5862,7295,9142,10113,10175,11822,12577,13055,15575,15935,
27,511,1536,1959,2959,4416,5040,5863,7296,9143,10114,10176,11823,12578,13056,15576,15936,
28,512,1537,1960,2960,4417,5041,5864,7297,9144,10115,10177,11824,12579,13057,15577,15937,
29,513,1538,1961,2961,4418,5042,5865,7298,9145,10116,10178,11825,12580,13058,15578,15938,
30,514,1539,1962,2962,4419,5043,5866,7299,9146,10117,10179,11826,12581,13059,15579,15939,
31,515,1540,1963,2963,4420,5044,5867,7300,9147,10118,10180,11827,12582,13060,15580,15940,
32,516,1541,1964,2964,4421,5045,5868,7301,9148,10119,10181,11828,12583,13061,15581,15941,
33,517,1542,1965,2965,4422,5046,5869,7302,9149,10120,10182,11829,12584,13062,15582,15942,
34,518,1543,1966,2966,4423,5047,5870,7303,9150,10121,10183,11830,12585,13063,15583,15943,
35,519,1544,1967,2967,4424,5048,5871,7304,9151,10122,10184,11831,12586,13064,15584,15944,
36,520,1545,1968,2968,4425,5049,5872,7305,9152,10123,10185,11832,12587,13065,15585,15945,
37,521,1546,1969,2969,4426,5050,5873,7306,9153,10124,10186,11833,12588,13066,15586,15946,
38,522,1547,1970,2970,4427,5051,5874,7307,9154,10125,10187,11834,12589,13067,15587,15947,
39,523,1548,1971,2971,4428,5052,5875,7308,9155,10126,10188,11835,12590,13068,15588,15948,
40,524,1549,1972,2972,4429,5053,5876,7309,9156,10127,10189,11836,12591,13069,15589,15949,
41,525,1550,1973,2973,4430,5054,5877,7310,9157,10128,10190,11837,12592,13070,15590,15950,
42,526,1551,1974,2974,4431,5055,5878,7311,9158,10129,10191,11838,12593,13071,15591,15951,
43,527,1552,1975,2975,4432,5056,5879,7312,9159,10130,10192,11839,12594,13072,15592,15952,
44,528,1553,1976,2976,4433,5057,5880,7313,9160,10131,10193,11840,12595,13073,15593,15953,
45,529,1554,1977,2977,4434,5058,5881,7314,9161,10132,10194,11841,12596,13074,15594,15954,
46,530,1555,1978,2978,4435,5059,5882,7315,9162,10133,10195,11842,12597,13075,15595,15955,
47,531,1556,1979,2979,4436,5060,5883,7316,9163,10134,10196,11843,12598,13076,15596,15956,
48,532,1557,1980,2980,4437,5061,5884,7317,9164,10135,10197,11844,12599,13077,15597,15957,
49,533,1558,1981,2981,4438,5062,5885,7318,9165,10136,10198,11845,12240,13078,15598,15958,
50,534,1559,1982,2982,4439,5063,5886,7319,9166,10137,10199,11846,12241,13079,15599,15959,
51,535,1560,1983,2983,4440,5064,5887,7320,9167,10138,10200,11847,12242,13080,15600,15960,
52,536,1561,1984,2984,4441,5065,5888,7321,9168,10139,10201,11848,12243,13081,15601,15961,
53,537,1562,1985,2985,4442,5066,5889,7322,9169,10140,10202,11849,12244,13082,15602,15962,
54,538,1563,1986,2986,4443,5067,5890,7323,9170,10141,10203,11850,12245,13083,15603,15963,
55,539,1564,1987,2987,4444,5068,5891,7324,9171,10142,10204,11851,12246,13084,15604,15964,
56,540,1565,1988,2988,4445,5069,5892,7325,9172,10143,10205,11852,12247,13085,15605,15965,
57,541,1566,1989,2989,4446,5070,5893,7326,9173,10144,10206,11853,12248,13086,15606,15966,
58,542,1567,1990,2990,4447,5071,5894,7327,9174,10145,10207,11854,12249,13087,15607,15967,
59,543,1568,1991,2991,4448,5072,5895,7328,9175,10146,10208,11855,12250,13088,15608,15968,
60,544,1569,1992,2992,4449,5073,5896,7329,9176,10147,10209,11856,12251,13089,15609,15969,
61,545,1570,1993,2993,4450,5074,5897,7330,9177,10148,10210,11857,12252,13090,15610,15970,
62,546,1571,1994,2994,4451,5075,5898,7331,9178,10149,10211,11858,12253,13091,15611,15971,
63,547,1572,1995,2995,4452,5076,5899,7332,9179,10150,10212,11859,12254,13092,15612,15972,
64,548,1573,1996,2996,4453,5077,5900,7333,9180,10151,10213,11860,12255,13093,15613,15973,
65,549,1574,1997,2997,4454,5078,5901,7334,9181,10152,10214,11861,12256,13094,15614,15974,
66,550,1575,1998,2998,4455,5079,5902,7335,9182,10153,10215,11862,12257,13095,15615,15975,
67,551,1576,1999,2999,4456,5080,5903,7336,9183,10154,10216,11863,12258,13096,15616,15976,
68,552,1577,2000,3000,4457,5081,5904,7337,9184,10155,10217,11864,12259,13097,15617,15977,
69,553,1578,2001,3001,4458,5082,5905,7338,9185,10156,10218,11865,12260,13098,15618,15978,
70,554,1579,2002,3002,4459,5083,5906,7339,9186,10157,10219,11866,12261,13099,15619,15979,
71,555,1580,2003,3003,4460,5084,5907,7340,9187,10158,10220,11867,12262,13100,15620,15980,
72,556,1581,2004,3004,4461,5085,5908,7341,9188,10159,10221,11868,12263,13101,15621,15981,
73,557,1582,2005,3005,4462,5086,5909,7342,9189,10160,10222,11869,12264,13102,15622,15982,
74,558,1583,2006,3006,4463,5087,5910,7343,9190,10161,10223,11870,12265,13103,15623,15983,
75,559,1584,2007,3007,4464,5088,5911,7344,9191,10162,10224,11871,12266,13104,15624,15984,
76,560,1585,2008,3008,4465,5089,5912,7345,9192,10163,10225,11872,12267,13105,15625,15985,
77,561,1586,2009,3009,4466,5090,5913,7346,9193,10164,10226,11873,12268,13106,15626,15986,
78,562,1587,2010,3010,4467,5091,5914,7347,9194,10165,10227,11874,12269,13107,15627,15987,
79,563,1588,2011,3011,4468,5092,5915,7348,9195,10166,10228,11875,12270,13108,15628,15988,
80,564,1589,2012,3012,4469,5093,5916,7349,9196,10167,10229,11876,12271,13109,15629,15989,
81,565,1590,2013,3013,4470,5094,5917,7350,9197,10168,10230,11877,12272,13110,15630,15990,
82,566,1591,2014,3014,4471,5095,5918,7351,9198,10169,10231,11878,12273,13111,15631,15991,
83,567,1592,2015,3015,4472,5096,5919,7352,9199,10170,10232,11879,12274,13112,15632,15992,
84,568,1593,2016,3016,4473,5097,5920,7353,9200,10171,10233,11520,12275,13113,15633,15993,
85,569,1594,2017,3017,4474,5098,5921,7354,9201,10172,10234,11521,12276,13114,15634,15994,
86,570,1595,2018,3018,4475,5099,5922,7355,9202,10173,10235,11522,12277,13115,15635,15995,
87,571,1596,2019,3019,4476,5100,5923,7356,9203,10174,10236,11523,12278,13116,15636,15996,
88,572,1597,2020,3020,4477,5101,5924,7357,9204,10175,10237,11524,12279,13117,15637,15997,
89,573,1598,2021,3021,4478,5102,5925,7358,9205,10176,10238,11525,12280,13118,15638,15998,
90,574,1599,2022,3022,4479,5103,5926,7359,9206,10177,10239,11526,12281,13119,15639,15999,
91,575,1600,2023,3023,4480,5104,5927,7360,9207,10178,10240,11527,12282,13120,15640,16000,
92,576,1601,2024,3024,4481,5105,5928,7361,9208,10179,10241,11528,12283,13121,15641,16001,
93,577,1602,2025,3025,4482,5106,5929,7362,9209,10180,10242,11529,12284,13122,15642,16002,
94,578,1603,2026,3026,4483,5107,5930,7363,9210,10181,10243,11530,12285,13123,15643,16003,
95,579,1604,2027,3027,4484,5108,5931,7364,9211,10182,10244,11531,12286,13124,15644,16004,
96,580,1605,2028,3028,4485,5109,5932,7365,9212,10183,10245,11532,12287,13125,15645,16005,
97,581,1606,2029,3029,4486,5110,5933,7366,9213,10184,10246,11533,12288,13126,15646,16006,
98,582,1607,2030,3030,4487,5111,5934,7367,9214,10185,10247,11534,12289,13127,15647,16007,
99,583,1608,2031,3031,4488,5112,5935,7368,9215,10186,10248,11535,12290,13128,15648,16008,
100,584,1609,2032,3032,4489,5113,5936,7369,9216,10187,10249,11536,12291,13129,15649,16009,
101,585,1610,2033,3033,4490,5114,5937,7370,9217,10188,10250,11537,12292,13130,15650,16010,
102,586,1611,2034,3034,4491,5115,5938,7371,9218,10189,10251,11538,12293,13131,15651,16011,
103,587,1612,2035,3035,4492,5116,5939,7372,9219,10190,10252,11539,12294,13132,15652,16012,
104,588,1613,2036,3036,4493,5117,5940,7373,9220,10191,10253,11540,12295,13133,15653,16013,
105,589,1614,2037,3037,4494,5118,5941,7374,9221,10192,10254,11541,12296,13134,15654,16014,
106,590,1615,2038,3038,4495,5119,5942,7375,9222,10193,10255,11542,12297,13135,15655,16015,
107,591,1616,2039,3039,4496,5120,5943,7376,9223,10194,10256,11543,12298,13136,15656,16016,
108,592,1617,2040,3040,4497,5121,5944,7377,9224,10195,10257,11544,12299,13137,15657,16017,
109,593,1618,2041,3041,4498,5122,5945,7378,9225,10196,10258,11545,12300,13138,15658,16018,
110,594,1619,2042,3042,4499,5123,5946,7379,9226,10197,10259,11546,12301,13139,15659,16019,
111,595,1620,2043,3043,4500,5124,5947,7380,9227,10198,10260,11547,12302,13140,15660,16020,
112,596,1621,2044,3044,4501,5125,5948,7381,9228,10199,10261,11548,12303,13141,15661,16021,
113,597,1622,2045,3045,4502,5126,5949,7382,9229,10200,10262,11549,12304,13142,15662,16022,
114,598,1623,2046,3046,4503,5127,5950,7383,9230,10201,10263,11550,12305,13143,15663,16023,
115,599,1624,2047,3047,4504,5128,5951,7384,9231,10202,10264,11551,12306,13144,15664,16024,
116,600,1625,2048,3048,4505,5129,5952,7385,9232,10203,10265,11552,12307,13145,15665,16025,
117,601,1626,2049,3049,4506,5130,5953,7386,9233,10204,10266,11553,12308,13146,15666,16026,
118,602,1627,2050,3050,4507,5131,5954,7387,9234,10205,10267,11554,12309,13147,15667,16027,
119,603,1628,2051,3051,4508,5132,5955,7388,9235,10206,10268,11555,12310,13148,15668,16028,
120,604,1629,2052,3052,4509,5133,5956,7389,9236,10207,10269,11556,12311,13149,15669,16029,
121,605,1630,2053,3053,4510,5134,5957,7390,9237,10208,10270,11557,12312,13150,15670,16030,
122,606,1631,2054,3054,4511,5135,5958,7391,9238,10209,10271,11558,12313,13151,15671,16031,
123,607,1632,2055,3055,4512,5136,5959,7392,9239,10210,10272,11559,12314,13152,15672,16032,
124,608,1633,2056,3056,4513,5137,5960,7393,9240,10211,10273,11560,12315,13153,15673,16033,
125,609,1634,2057,3057,4514,5138,5961,7394,9241,10212,10274,11561,12316,13154,15674,16034,
126,610,1635,2058,3058,4515,5139,5962,7395,9242,10213,10275,11562,12317,13155,15675,16035,
127,611,1636,2059,3059,4516,5140,5963,7396,9243,10214,10276,11563,12318,13156,15676,16036,
128,612,1637,2060,3060,4517,5141,5964,7397,9244,10215,10277,11564,12319,13157,15677,16037,
129,613,1638,2061,3061,4518,5142,5965,7398,9245,10216,10278,11565,12320,13158,15678,16038,
130,614,1639,2062,3062,4519,5143,5966,7399,9246,10217,10279,11566,12321,13159,15679,16039,
131,615,1640,2063,3063,4520,5144,5967,7400,9247,10218,10280,11567,12322,13160,15680,16040,
132,616,1641,2064,3064,4521,5145,5968,7401,9248,10219,10281,11568,12323,13161,15681,16041,
133,617,1642,2065,3065,4522,5146,5969,7402,9249,10220,10282,11569,12324,13162,15682,16042,
134,618,1643,2066,3066,4523,5147,5970,7403,9250,10221,10283,11570,12325,13163,15683,16043,
135,619,1644,2067,3067,4524,5148,5971,7404,9251,10222,10284,11571,12326,13164,15684,16044,
136,620,1645,2068,3068,4525,5149,5972,7405,9252,10223,10285,11572,12327,13165,15685,16045,
137,621,1646,2069,3069,4526,5150,5973,7406,9253,10224,10286,11573,12328,13166,15686,16046,
138,622,1647,2070,3070,4527,5151,5974,7407,9254,10225,10287,11574,12329,13167,15687,16047,
139,623,1648,2071,3071,4528,5152,5975,7408,9255,10226,10288,11575,12330,13168,15688,16048,
140,624,1649,2072,3072,4529,5153,5976,7409,9256,10227,10289,11576,12331,13169,15689,16049,
141,625,1650,2073,3073,4530,5154,5977,7410,9257,10228,10290,11577,12332,13170,15690,16050,
142,626,1651,2074,3074,4531,5155,5978,7411,9258,10229,10291,11578,12333,13171,15691,16051,
143,627,1652,2075,3075,4532,5156,5979,7412,9259,10230,10292,11579,12334,13172,15692,16052,
144,628,1653,2076,3076,4533,5157,5980,7413,9260,10231,10293,11580,12335,13173,15693,16053,
145,629,1654,2077,3077,4534,5158,5981,7414,9261,10232,10294,11581,12336,13174,15694,16054,
146,630,1655,2078,3078,4535,5159,5982,7415,9262,10233,10295,11582,12337,13175,15695,16055,
147,631,1656,2079,3079,4536,5160,5983,7416,9263,10234,10296,11583,12338,13176,15696,16056,
148,632,1657,2080,3080,4537,5161,5984,7417,9264,10235,10297,11584,12339,13177,15697,16057,
149,633,1658,2081,3081,4538,5162,5985,7418,9265,10236,10298,11585,12340,13178,15698,16058,
150,634,1659,2082,3082,4539,5163,5986,7419,9266,10237,10299,11586,12341,13179,15699,16059,
151,635,1660,2083,3083,4540,5164,5987,7420,9267,10238,10300,11587,12342,13180,15700,16060,
152,636,1661,2084,3084,4541,5165,5988,7421,9268,10239,10301,11588,12343,13181,15701,16061,
153,637,1662,2085,3085,4542,5166,5989,7422,9269,10240,10302,11589,12344,13182,15702,16062,
154,638,1663,2086,3086,4543,5167,5990,7423,9270,10241,10303,11590,12345,13183,15703,16063,
155,639,1664,2087,3087,4544,5168,5991,7424,9271,10242,10304,11591,12346,13184,15704,16064,
156,640,1665,2088,3088,4545,5169,5992,7425,9272,10243,10305,11592,12347,13185,15705,16065,
157,641,1666,2089,3089,4546,5170,5993,7426,9273,10244,10306,11593,12348,13186,15706,16066,
158,642,1667,2090,3090,4547,5171,5994,7427,9274,10245,10307,11594,12349,13187,15707,16067,
159,643,1668,2091,3091,4548,5172,5995,7428,9275,10246,10308,11595,12350,13188,15708,16068,
160,644,1669,2092,3092,4549,5173,5996,7429,9276,10247,10309,11596,12351,13189,15709,16069,
161,645,1670,2093,3093,4550,5174,5997,7430,9277,10248,10310,11597,12352,13190,15710,16070,
162,646,1671,2094,3094,4551,5175,5998,7431,9278,10249,10311,11598,12353,13191,15711,16071,
163,647,1672,2095,3095,4552,5176,5999,7432,9279,10250,10312,11599,12354,13192,15712,16072,
164,648,1673,2096,3096,4553,5177,6000,7433,9280,10251,10313,11600,12355,13193,15713,16073,
165,649,1674,2097,3097,4554,5178,6001,7434,9281,10252,10314,11601,12356,13194,15714,16074,
166,650,1675,2098,3098,4555,5179,6002,7435,9282,10253,10315,11602,12357,13195,15715,16075,
167,651,1676,2099,3099,4556,5180,6003,7436,9283,10254,10316,11603,12358,13196,15716,16076,
168,652,1677,2100,3100,4557,5181,6004,7437,9284,10255,10317,11604,12359,13197,15717,16077,
169,653,1678,2101,3101,4558,5182,6005,7438,9285,10256,10318,11605,12360,13198,15718,16078,
170,654,1679,2102,3102,4559,5183,6006,7439,9286,10257,10319,11606,12361,13199,15719,16079,
171,655,1680,2103,3103,4560,5184,6007,7440,9287,10258,10320,11607,12362,13200,15720,16080,
172,656,1681,2104,3104,4561,5185,6008,7441,9288,10259,10321,11608,12363,13201,15721,16081,
173,657,1682,2105,3105,4562,5186,6009,7442,9289,10260,10322,11609,12364,13202,15722,16082,
174,658,1683,2106,3106,4563,5187,6010,7443,9290,10261,10323,11610,12365,13203,15723,16083,
175,659,1684,2107,3107,4564,5188,6011,7444,9291,10262,10324,11611,12366,13204,15724,16084,
176,660,1685,2108,3108,4565,5189,6012,7445,9292,10263,10325,11612,12367,13205,15725,16085,
177,661,1686,2109,3109,4566,5190,6013,7446,9293,10264,10326,11613,12368,13206,15726,16086,
178,662,1687,2110,3110,4567,5191,6014,7447,9294,10265,10327,11614,12369,13207,15727,16087,
179,663,1688,2111,3111,4568,5192,6015,7448,9295,10266,10328,11615,12370,13208,15728,16088,
180,664,1689,2112,3112,4569,5193,6016,7449,9296,10267,10329,11616,12371,13209,15729,16089,
181,665,1690,2113,3113,4570,5194,6017,7450,9297,10268,10330,11617,12372,13210,15730,16090,
182,666,1691,2114,3114,4571,5195,6018,7451,9298,10269,10331,11618,12373,13211,15731,16091,
183,667,1692,2115,3115,4572,5196,6019,7452,9299,10270,10332,11619,12374,13212,15732,16092,
184,668,1693,2116,3116,4573,5197,6020,7453,9300,10271,10333,11620,12375,13213,15733,16093,
185,669,1694,2117,3117,4574,5198,6021,7454,9301,10272,10334,11621,12376,13214,15734,16094,
186,670,1695,2118,3118,4575,5199,6022,7455,9302,10273,10335,11622,12377,13215,15735,16095,
187,671,1696,2119,3119,4576,5200,6023,7456,9303,10274,10336,11623,12378,13216,15736,16096,
188,672,1697,2120,3120,4577,5201,6024,7457,9304,10275,10337,11624,12379,13217,15737,16097,
189,673,1698,2121,3121,4578,5202,6025,7458,9305,10276,10338,11625,12380,13218,15738,16098,
190,674,1699,2122,3122,4579,5203,6026,7459,9306,10277,10339,11626,12381,13219,15739,16099,
191,675,1700,2123,3123,4580,5204,6027,7460,9307,10278,10340,11627,12382,13220,15740,16100,
192,676,1701,2124,3124,4581,5205,6028,7461,9308,10279,10341,11628,12383,13221,15741,16101,
193,677,1702,2125,3125,4582,5206,6029,7462,9309,10280,10342,11629,12384,13222,15742,16102,
194,678,1703,2126,3126,4583,5207,6030,7463,9310,10281,10343,11630,12385,13223,15743,16103,
195,679,1704,2127,3127,4584,5208,6031,7464,9311,10282,10344,11631,12386,13224,15744,16104,
196,680,1705,2128,3128,4585,5209,6032,7465,9312,10283,10345,11632,12387,13225,15745,16105,
197,681,1706,2129,3129,4586,5210,6033,7466,9313,10284,10346,11633,12388,13226,15746,16106,
198,682,1707,2130,3130,4587,5211,6034,7467,9314,10285,10347,11634,12389,13227,15747,16107,
199,683,1708,2131,3131,4588,5212,6035,7468,9315,10286,10348,11635,12390,13228,15748,16108,
200,684,1709,2132,3132,4589,5213,6036,7469,9316,10287,10349,11636,12391,13229,15749,16109,
201,685,1710,2133,3133,4590,5214,6037,7470,9317,10288,10350,11637,12392,13230,15750,16110,
202,686,1711,2134,3134,4591,5215,6038,7471,9318,10289,10351,11638,12393,13231,15751,16111,
203,687,1712,2135,3135,4592,5216,6039,7472,9319,10290,10352,11639,12394,13232,15752,16112,
204,688,1713,2136,3136,4593,5217,6040,7473,9320,10291,10353,11640,12395,13233,15753,16113,
205,689,1714,2137,3137,4594,5218,6041,7474,9321,10292,10354,11641,12396,13234,15754,16114,
206,690,1715,2138,3138,4595,5219,6042,7475,9322,10293,10355,11642,12397,13235,15755,16115,
207,691,1716,2139,3139,4596,5220,6043,7476,9323,10294,10356,11643,12398,13236,15756,16116,
208,692,1717,2140,3140,4597,5221,6044,7477,9324,10295,10357,11644,12399,13237,15757,16117,
209,693,1718,2141,3141,4598,5222,6045,7478,9325,10296,10358,11645,12400,13238,15758,16118,
210,694,1719,2142,3142,4599,5223,6046,7479,9326,10297,10359,11646,12401,13239,15759,16119,
211,695,1720,2143,3143,4600,5224,6047,7480,9327,10298,10360,11647,12402,13240,15760,16120,
212,696,1721,2144,3144,4601,5225,6048,7481,9328,10299,10361,11648,12403,13241,15761,16121,
213,697,1722,2145,3145,4602,5226,6049,7482,9329,10300,10362,11649,12404,13242,15762,16122,
214,698,1723,2146,3146,4603,5227,6050,7483,9330,10301,10363,11650,12405,13243,15763,16123,
215,699,1724,2147,3147,4604,5228,6051,7484,9331,10302,10364,11651,12406,13244,15764,16124,
216,700,1725,2148,3148,4605,5229,6052,7485,9332,10303,10365,11652,12407,13245,15765,16125,
217,701,1726,2149,3149,4606,5230,6053,7486,9333,10304,10366,11653,12408,13246,15766,16126,
218,702,1727,2150,3150,4607,5231,6054,7487,9334,10305,10367,11654,12409,13247,15767,16127,
219,703,1728,2151,3151,4608,5232,6055,7488,9335,10306,10368,11655,12410,13248,15768,16128,
220,704,1729,2152,3152,4609,5233,6056,7489,9336,10307,10369,11656,12411,13249,15769,16129,
221,705,1730,2153,3153,4610,5234,6057,7490,9337,10308,10370,11657,12412,13250,15770,16130,
222,706,1731,2154,3154,4611,5235,6058,7491,9338,10309,10371,11658,12413,13251,15771,16131,
223,707,1732,2155,3155,4612,5236,6059,7492,9339,10310,10372,11659,12414,13252,15772,16132,
224,708,1733,2156,3156,4613,5237,6060,7493,9340,10311,10373,11660,12415,13253,15773,16133,
225,709,1734,2157,3157,4614,5238,6061,7494,9341,10312,10374,11661,12416,13254,15774,16134,
226,710,1735,2158,3158,4615,5239,6062,7495,9342,10313,10375,11662,12417,13255,15775,16135,
227,711,1736,2159,3159,4616,5240,6063,7496,9343,10314,10376,11663,12418,13256,15776,16136,
228,712,1737,1800,3160,4617,5241,6064,7497,9344,10315,10377,11664,12419,13257,15777,16137,
229,713,1738,1801,3161,4618,5242,6065,7498,9345,10316,10378,11665,12420,13258,15778,16138,
230,714,1739,1802,3162,4619,5243,6066,7499,9346,10317,10379,11666,12421,13259,15779,16139,
231,715,1740,1803,3163,4620,5244,6067,7500,9347,10318,10380,11667,12422,13260,15780,16140,
232,716,1741,1804,3164,4621,5245,6068,7501,9348,10319,10381,11668,12423,13261,15781,16141,
233,717,1742,1805,3165,4622,5246,6069,7502,9349,10320,10382,11669,12424,13262,15782,16142,
234,718,1743,1806,3166,4623,5247,6070,7503,9350,10321,10383,11670,12425,13263,15783,16143,
235,719,1744,1807,3167,4624,5248,6071,7504,9351,10322,10384,11671,12426,13264,15784,16144,
236,360,1745,1808,3168,4625,5249,6072,7505,9352,10323,10385,11672,12427,13265,15785,16145,
237,361,1746,1809,3169,4626,5250,6073,7506,9353,10324,10386,11673,12428,13266,15786,16146,
238,362,1747,1810,3170,4627,5251,6074,7507,9354,10325,10387,11674,12429,13267,15787,16147,
239,363,1748,1811,3171,4628,5252,6075,7508,9355,10326,10388,11675,12430,13268,15788,16148,
240,364,1749,1812,3172,4629,5253,6076,7509,9356,10327,10389,11676,12431,13269,15789,16149,
241,365,1750,1813,3173,4630,5254,6077,7510,9357,10328,10390,11677,12432,13270,15790,16150,
242,366,1751,1814,3174,4631,5255,6078,7511,9358,10329,10391,11678,12433,13271,15791,16151,
243,367,1752,1815,3175,4632,5256,6079,7512,9359,10330,10392,11679,12434,13272,15792,16152,
244,368,1753,1816,3176,4633,5257,6080,7513,9000,10331,10393,11680,12435,13273,15793,16153,
245,369,1754,1817,3177,4634,5258,6081,7514,9001,10332,10394,11681,12436,13274,15794,16154,
246,370,1755,1818,3178,4635,5259,6082,7515,9002,10333,10395,11682,12437,13275,15795,16155,
247,371,1756,1819,3179,4636,5260,6083,7516,9003,10334,10396,11683,12438,13276,15796,16156,
248,372,1757,1820,3180,4637,5261,6084,7517,9004,10335,10397,11684,12439,13277,15797,16157,
249,373,1758,1821,3181,4638,5262,6085,7518,9005,10336,10398,11685,12440,13278,15798,16158,
250,374,1759,1822,3182,4639,5263,6086,7519,9006,10337,10399,11686,12441,13279,15799,16159,
251,375,1760,1823,3183,4640,5264,6087,7520,9007,10338,10400,11687,12442,13280,15800,16160,
252,376,1761,1824,3184,4641,5265,6088,7521,9008,10339,10401,11688,12443,13281,15801,16161,
253,377,1762,1825,3185,4642,5266,6089,7522,9009,10340,10402,11689,12444,13282,15802,16162,
254,378,1763,1826,3186,4643,5267,6090,7523,9010,10341,10403,11690,12445,13283,15803,16163,
255,379,1764,1827,3187,4644,5268,6091,7524,9011,10342,10404,11691,12446,13284,15804,16164,
256,380,1765,1828,3188,4645,5269,6092,7525,9012,10343,10405,11692,12447,13285,15805,16165,
257,381,1766,1829,3189,4646,5270,6093,7526,9013,10344,10406,11693,12448,13286,15806,16166,
258,382,1767,1830,3190,4647,5271,6094,7527,9014,10345,10407,11694,12449,13287,15807,16167,
259,383,1768,1831,3191,4648,5272,6095,7528,9015,10346,10408,11695,12450,13288,15808,16168,
260,384,1769,1832,3192,4649,5273,6096,7529,9016,10347,10409,11696,12451,13289,15809,16169,
261,385,1770,1833,3193,4650,5274,6097,7530,9017,10348,10410,11697,12452,13290,15810,16170,
262,386,1771,1834,3194,4651,5275,6098,7531,9018,10349,10411,11698,12453,13291,15811,16171,
263,387,1772,1835,3195,4652,5276,6099,7532,9019,10350,10412,11699,12454,13292,15812,16172,
264,388,1773,1836,3196,4653,5277,6100,7533,9020,10351,10413,11700,12455,13293,15813,16173,
265,389,1774,1837,3197,4654,5278,6101,7534,9021,10352,10414,11701,12456,13294,15814,16174,
266,390,1775,1838,3198,4655,5279,6102,7535,9022,10353,10415,11702,12457,13295,15815,16175,
267,391,1776,1839,3199,4656,5280,6103,7536,9023,10354,10416,11703,12458,13296,15816,16176,
268,392,1777,1840,3200,4657,5281,6104,7537,9024,10355,10417,11704,12459,13297,15817,16177,
269,393,1778,1841,3201,4658,5282,6105,7538,9025,10356,10418,11705,12460,13298,15818,16178,
270,394,1779,1842,3202,4659,5283,6106,7539,9026,10357,10419,11706,12461,13299,15819,16179,
271,395,1780,1843,3203,4660,5284,6107,7540,9027,10358,10420,11707,12462,13300,15820,16180,
272,396,1781,1844,3204,4661,5285,6108,7541,9028,10359,10421,11708,12463,13301,15821,16181,
273,397,1782,1845,3205,4662,5286,6109,7542,9029,10360,10422,11709,12464,13302,15822,16182,
274,398,1783,1846,3206,4663,5287,6110,7543,9030,10361,10423,11710,12465,13303,15823,16183,
275,399,1784,1847,3207,4664,5288,6111,7544,9031,10362,10424,11711,12466,13304,15824,16184,
276,400,1785,1848,3208,4665,5289,6112,7545,9032,10363,10425,11712,12467,13305,15825,16185,
277,401,1786,1849,3209,4666,5290,6113,7546,9033,10364,10426,11713,12468,13306,15826,16186,
278,402,1787,1850,3210,4667,5291,6114,7547,9034,10365,10427,11714,12469,13307,15827,16187,
279,403,1788,1851,3211,4668,5292,6115,7548,9035,10366,10428,11715,12470,13308,15828,16188,
280,404,1789,1852,3212,4669,5293,6116,7549,9036,10367,10429,11716,12471,13309,15829,16189,
281,405,1790,1853,3213,4670,5294,6117,7550,9037,10368,10430,11717,12472,13310,15830,16190,
282,406,1791,1854,3214,4671,5295,6118,7551,9038,10369,10431,11718,12473,13311,15831,16191,
283,407,1792,1855,3215,4672,5296,6119,7552,9039,10370,10432,11719,12474,13312,15832,16192,
284,408,1793,1856,3216,4673,5297,5760,7553,9040,10371,10433,11720,12475,13313,15833,16193,
285,409,1794,1857,3217,4674,5298,5761,7554,9041,10372,10434,11721,12476,13314,15834,16194,
286,410,1795,1858,3218,4675,5299,5762,7555,9042,10373,10435,11722,12477,13315,15835,16195,
287,411,1796,1859,3219,4676,5300,5763,7556,9043,10374,10436,11723,12478,13316,15836,16196,
288,412,1797,1860,3220,4677,5301,5764,7557,9044,10375,10437,11724,12479,13317,15837,16197,
289,413,1798,1861,3221,4678,5302,5765,7558,9045,10376,10438,11725,12480,13318,15838,16198,
290,414,1799,1862,3222,4679,5303,5766,7559,9046,10377,10439,11726,12481,13319,15839,16199,
		others => 0);
	end function;
end package body;
