-- code table generated from table_vector.txt by generate_table_vector_vhd.cc
--
-- Copyright 2019 Ahmet Inan <inan@aicodix.de>

use work.ldpc_scalar.all;
use work.ldpc_vector.all;

package table_vector is
	function init_vector_parities return vector_parities;
	function init_vector_counts return vector_counts;
	function init_vector_offsets return vector_offsets;
	function init_vector_shifts return vector_shifts;
end package;

package body table_vector is
	function init_vector_parities return vector_parities is
	begin
		return 135;
	end function;

	function init_vector_counts return vector_counts is
	begin
		return (
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
14,
		others => count_scalar'low);
	end function;

	function init_vector_offsets return vector_offsets is
	begin
		return (
3,7,13,33,123,131,218,223,266,345,346,401,533,536,
5,28,37,40,43,111,164,230,246,304,381,399,513,516,
12,24,26,31,38,64,159,165,267,288,294,349,426,429,
4,22,36,47,131,134,182,225,269,279,395,404,536,539,
1,17,18,69,70,108,167,194,204,318,327,339,471,474,
3,29,38,41,44,112,162,228,247,305,382,400,514,517,
14,23,30,47,56,79,182,205,258,307,317,375,449,452,
0,15,25,33,46,69,168,169,171,291,303,367,435,438,
5,6,12,35,125,130,217,222,265,345,347,400,532,535,
14,30,34,40,40,124,159,175,205,310,321,330,442,445,
18,24,29,62,81,104,142,216,221,293,351,354,483,486,
15,16,17,28,91,97,150,220,232,284,285,393,417,420,
5,6,9,25,52,96,137,211,231,359,366,382,498,501,
3,21,38,46,130,133,181,227,268,281,394,403,535,538,
17,20,26,29,36,49,145,155,269,290,294,319,422,425,
8,10,11,53,86,117,188,207,265,306,323,388,455,458,
30,43,43,99,111,126,157,197,234,285,369,391,501,504,
3,6,13,19,28,88,163,172,263,298,324,335,430,433,
4,7,14,34,48,63,168,198,248,311,331,333,465,468,
1,2,33,38,40,121,183,201,256,309,363,391,523,526,
3,9,21,29,117,122,138,188,247,273,341,387,405,408,
11,18,18,30,60,90,197,210,225,275,360,379,492,495,
16,19,25,28,38,48,144,154,268,289,296,318,421,424,
5,23,37,45,129,132,180,226,267,280,393,402,534,537,
4,8,11,24,51,98,136,210,233,358,368,381,500,503,
7,9,10,52,85,119,187,209,264,308,322,387,454,457,
15,16,17,27,90,96,152,219,231,283,287,395,419,422,
4,14,29,32,38,39,167,189,234,298,301,302,434,437,
12,31,35,41,41,125,160,176,206,311,322,331,443,446,
19,20,23,34,43,55,151,180,190,325,359,364,457,460,
0,21,42,42,77,79,174,201,214,349,362,386,481,484,
2,6,13,25,29,68,203,245,252,296,338,360,470,473,
8,14,31,33,87,108,136,139,149,284,300,323,416,419,
1,16,26,34,47,70,169,170,172,292,304,368,436,439,
21,28,39,44,59,99,141,156,198,291,324,370,423,426,
13,24,25,32,36,65,160,166,268,289,295,350,427,430,
2,15,34,37,55,87,147,222,242,278,313,357,489,492,
31,42,44,77,85,129,215,220,226,338,355,386,487,490,
3,6,8,22,92,121,141,154,255,272,276,343,408,411,
0,7,14,26,27,66,201,243,253,294,336,361,468,471,
16,24,31,61,81,115,140,196,222,331,341,397,463,466,
1,22,43,43,75,80,175,202,215,350,360,384,482,485,
3,12,37,41,57,107,192,231,262,290,327,381,459,462,
4,7,14,20,29,89,164,173,261,299,325,333,431,434,
10,18,18,27,49,106,184,253,257,274,319,344,451,454,
6,9,11,51,84,118,186,208,266,307,321,389,453,456,
4,13,38,39,58,105,193,232,263,288,328,382,460,463,
5,7,8,21,91,120,143,153,257,271,278,342,410,413,
1,22,32,57,97,119,148,249,254,304,333,389,521,524,
23,30,43,64,100,115,192,250,265,376,385,390,517,520,
19,25,27,60,82,102,143,217,219,291,352,355,484,487,
26,28,34,67,77,128,212,238,245,276,347,354,479,482,
5,14,36,40,59,106,194,233,261,289,329,383,461,464,
0,7,10,19,32,95,135,179,208,270,283,378,405,539,
25,27,33,66,76,127,211,237,244,278,346,356,478,481,
5,11,23,28,119,121,140,187,246,275,340,389,407,410,
22,32,42,63,99,114,194,249,264,375,384,392,516,519,
30,43,44,76,84,131,214,219,225,337,354,385,486,489,
5,8,12,35,49,64,169,199,246,309,332,334,466,469,
0,2,34,36,41,122,184,202,257,310,364,392,524,527,
3,7,10,26,53,97,135,212,232,357,367,383,499,502,
13,22,32,46,55,78,181,204,260,306,316,377,448,451,
16,24,34,40,123,133,218,249,258,287,393,398,525,528,
9,19,19,31,61,91,195,211,226,273,361,380,493,496,
10,15,18,39,85,109,198,239,244,353,372,379,511,514,
4,8,14,34,124,129,216,224,264,346,347,399,531,534,
21,31,44,65,101,116,193,251,266,377,386,391,518,521,
9,17,20,41,84,108,200,238,243,352,374,378,510,513,
4,6,7,23,90,122,142,155,256,270,277,344,409,412,
0,1,35,37,39,120,185,203,255,311,365,390,522,525,
3,5,10,73,73,126,163,189,261,281,353,396,528,531,
9,15,34,44,80,107,159,242,258,337,367,377,509,512,
17,25,32,62,82,116,138,197,223,332,339,398,464,467,
2,23,30,58,98,117,149,250,252,305,334,387,519,522,
6,22,36,103,103,113,174,185,238,317,327,373,505,508,
4,5,9,72,72,128,162,191,263,280,352,398,530,533,
1,8,11,20,30,93,136,177,209,271,284,379,406,537,
0,21,31,59,96,118,147,251,253,303,335,388,520,523,
15,16,17,29,92,98,151,221,233,282,286,394,418,421,
5,12,27,30,36,40,165,190,235,299,300,302,432,435,
20,26,28,61,83,103,141,218,220,292,353,356,485,488,
17,25,35,41,124,134,216,250,259,285,394,396,526,529,
2,23,44,44,76,78,176,203,213,348,361,385,480,483,
11,16,19,40,86,110,199,237,245,351,373,380,512,515,
0,6,36,38,41,93,157,171,228,271,306,312,438,441,
15,18,24,27,37,50,146,153,267,288,295,320,420,423,
1,14,23,40,94,134,177,213,229,298,364,402,496,499,
10,12,38,41,44,66,155,179,187,314,317,349,446,449,
0,27,35,72,82,116,207,235,240,342,372,401,474,477,
7,23,37,104,104,111,175,183,239,315,328,374,506,509,
1,17,33,36,54,89,149,224,241,277,312,359,491,494,
11,19,19,28,50,107,185,254,255,275,320,342,452,455,
31,44,44,100,112,127,158,195,235,286,370,392,502,505,
13,32,33,39,39,123,161,174,204,309,323,332,441,444,
10,16,35,42,78,105,160,240,259,338,368,375,507,510,
1,8,12,24,28,67,202,244,254,295,337,362,469,472,
2,6,9,18,31,94,137,178,207,272,282,380,407,538,
11,17,33,43,79,106,161,241,260,336,366,376,508,511,
4,27,36,39,42,113,163,229,248,303,383,401,515,518,
6,12,32,34,88,109,137,140,147,282,301,321,414,417,
7,13,30,35,89,110,135,138,148,283,302,322,415,418,
8,21,38,102,102,112,176,184,237,316,329,372,504,507,
11,15,22,26,26,53,145,146,150,281,371,403,413,416,
10,20,20,32,62,92,196,212,227,274,362,378,494,497,
3,6,13,33,50,65,170,200,247,310,330,335,467,470,
14,25,26,30,37,63,161,167,269,290,296,348,428,431,
2,12,21,41,95,132,178,214,230,299,365,403,497,500,
0,16,35,38,56,88,148,223,240,276,314,358,490,493,
4,10,22,27,118,120,139,186,248,274,339,388,406,409,
2,15,19,70,71,109,165,192,205,319,328,340,472,475,
9,16,23,24,24,51,144,146,151,279,369,404,411,414,
11,13,36,39,42,67,153,177,188,312,315,350,444,447,
1,28,33,73,83,114,208,236,241,343,373,399,475,478,
23,27,41,43,58,101,143,158,200,293,326,369,425,428,
2,8,37,38,40,95,156,173,230,270,308,314,440,443,
18,19,22,33,42,54,150,182,189,324,358,363,456,459,
24,29,35,68,75,126,210,239,243,277,345,355,477,480,
0,16,20,69,71,110,166,193,206,320,329,341,473,476,
5,8,12,18,27,87,162,171,262,297,326,334,429,432,
1,7,36,37,39,94,158,172,229,272,307,313,439,442,
2,29,34,74,81,115,209,234,242,344,374,400,476,479,
32,42,42,101,113,128,156,196,236,287,371,390,503,506,
10,17,21,25,25,52,144,145,152,280,370,402,412,415,
9,20,20,29,48,105,183,252,256,273,318,343,450,453,
32,42,43,75,86,130,213,221,227,336,356,384,488,491,
0,13,22,39,93,133,179,215,228,297,363,404,495,498,
15,26,30,60,83,114,139,195,224,330,340,396,462,465,
2,17,24,35,45,71,168,170,173,293,305,366,437,440,
3,13,28,31,37,41,166,191,236,297,300,301,433,436,
15,26,33,39,125,132,217,251,260,286,395,397,527,530,
22,29,40,42,57,100,142,157,199,292,325,371,424,427,
18,20,21,35,44,56,152,181,191,326,357,365,458,461,
3,4,11,74,74,127,164,190,262,279,351,397,529,532,
9,14,37,40,43,68,154,178,186,313,316,348,445,448,
12,21,31,45,54,80,180,206,259,308,315,376,447,450,
		others => 0);
	end function;

	function init_vector_shifts return vector_shifts is
	begin
		return (
101,108,105,65,87,0,34,16,0,10,55,0,0,0,
25,96,100,61,84,0,9,16,0,36,0,82,0,0,
108,0,93,45,10,87,0,107,63,63,0,71,0,0,
67,116,83,97,62,0,64,50,0,108,75,0,0,0,
81,65,62,0,53,112,5,57,0,91,28,0,0,0,
26,96,100,61,84,0,10,17,0,36,0,82,0,0,
111,31,72,0,13,75,0,77,7,94,0,102,0,0,
114,80,77,0,31,64,0,107,28,101,0,29,0,0,
100,108,105,64,86,0,34,16,0,55,9,0,0,0,
51,52,106,0,54,37,83,0,107,0,86,27,0,0,
61,15,83,95,0,22,59,0,63,61,0,118,0,0,
0,27,109,66,94,18,0,1,30,109,0,8,0,0,
35,62,92,94,21,0,112,73,0,70,0,69,0,0,
67,116,82,97,62,0,64,49,0,107,75,0,0,0,
15,0,52,116,56,21,97,0,74,0,85,100,0,0,
8,22,14,0,56,64,0,10,103,37,0,45,0,0,
45,8,37,0,105,74,30,110,0,52,0,84,0,0,
18,73,40,90,0,25,0,116,111,0,30,90,0,0,
105,73,63,38,69,0,60,0,84,9,87,0,0,0,
73,37,42,67,92,0,74,91,0,101,14,0,0,0,
0,93,117,104,14,59,0,30,50,0,9,60,0,0,
108,76,95,65,91,0,15,79,0,17,0,72,0,0,
15,0,52,116,55,21,97,0,74,0,84,100,0,0,
66,115,82,97,62,0,64,49,0,107,75,0,0,0,
36,62,92,95,22,0,113,74,0,71,0,70,0,0,
8,22,14,0,56,63,0,9,103,36,0,45,0,0,
28,110,0,67,95,19,0,2,31,110,0,8,0,0,
7,84,71,0,93,117,0,61,6,32,107,0,0,0,
52,52,106,0,54,37,83,0,107,0,86,27,0,0,
44,43,52,40,13,0,16,48,0,0,17,35,0,0,
62,30,72,98,66,0,68,92,0,0,37,6,0,0,
100,20,36,76,66,0,0,59,100,4,0,33,0,0,
13,0,68,5,57,107,111,27,0,0,114,57,0,0,
114,80,77,0,31,64,0,107,28,101,0,29,0,0,
0,26,70,59,66,15,100,0,91,0,54,20,0,0,
108,94,0,45,11,87,0,107,63,63,0,71,0,0,
101,78,119,109,105,0,109,0,98,24,63,0,0,0,
67,4,55,67,0,57,88,0,23,57,0,16,0,0,
70,0,29,7,96,4,0,61,11,67,0,9,0,0,
100,19,35,75,66,0,0,59,99,4,0,32,0,0,
17,114,38,0,65,75,46,0,86,0,107,13,0,0,
62,30,72,98,67,0,68,92,0,0,38,7,0,0,
36,12,104,4,0,8,0,6,61,101,0,51,0,0,
18,73,40,90,0,25,0,116,112,0,30,91,0,0,
66,55,86,48,0,81,0,57,57,91,0,67,0,0,
8,14,21,0,56,63,0,9,102,36,0,44,0,0,
36,12,104,5,0,9,0,6,61,102,0,51,0,0,
70,30,0,8,97,5,0,62,11,68,0,10,0,0,
66,105,23,89,76,0,118,85,0,52,111,0,0,0,
26,117,19,74,39,0,99,0,56,37,0,32,0,0,
61,15,84,96,0,23,59,0,64,62,0,118,0,0,
74,85,35,17,0,19,0,7,98,64,0,26,0,0,
36,12,105,5,0,9,0,6,62,102,0,51,0,0,
0,17,68,48,54,87,0,57,100,0,62,26,0,119,
74,85,35,17,0,19,0,7,98,63,0,25,0,0,
0,93,117,105,14,60,0,31,51,0,10,60,0,0,
26,116,19,74,39,0,98,0,56,37,0,31,0,0,
67,55,3,67,0,56,88,0,23,57,0,16,0,0,
105,73,64,38,69,0,60,0,85,10,87,0,0,0,
38,73,42,68,92,0,74,91,0,101,14,0,0,0,
36,62,92,94,21,0,113,73,0,71,0,69,0,0,
111,31,71,0,13,75,0,77,6,94,0,101,0,0,
50,58,61,114,0,33,29,38,0,76,0,60,0,0,
109,76,95,65,91,0,16,79,0,18,0,72,0,0,
62,3,7,59,102,0,18,65,0,117,13,0,0,0,
100,107,104,64,86,0,34,15,0,9,54,0,0,0,
27,117,19,74,39,0,99,0,56,37,0,32,0,0,
62,2,6,58,102,0,17,65,0,117,12,0,0,0,
70,30,0,7,97,4,0,61,11,68,0,9,0,0,
73,37,41,67,92,0,73,90,0,100,13,0,0,0,
114,117,55,15,98,0,26,53,0,59,83,0,0,0,
78,109,119,25,19,0,73,0,63,18,1,0,0,0,
17,114,38,0,65,75,47,0,86,0,108,13,0,0,
65,104,23,88,75,0,117,84,0,51,110,0,0,0,
21,65,3,0,102,112,90,36,0,23,78,0,0,0,
118,114,56,16,99,0,27,53,0,60,84,0,0,0,
0,17,68,48,55,88,0,58,100,0,62,26,0,0,
66,105,23,88,76,0,118,84,0,52,110,0,0,0,
110,0,27,66,94,18,0,1,30,110,0,8,0,0,
6,84,71,0,93,116,0,60,5,31,0,106,0,0,
61,15,84,96,0,23,60,0,64,62,0,118,0,0,
50,58,61,114,0,33,30,38,0,77,0,61,0,0,
61,29,71,97,66,0,67,91,0,0,37,6,0,0,
62,3,7,59,102,0,18,66,0,118,13,0,0,0,
96,61,0,83,100,17,8,0,49,94,0,62,0,0,
15,0,52,116,55,20,96,0,74,0,84,99,0,0,
12,7,87,89,0,100,110,27,0,43,0,13,0,0,
33,49,2,22,0,101,1,0,110,0,75,57,0,0,
21,95,10,0,12,48,0,55,5,0,23,37,0,0,
21,65,3,0,102,113,90,37,0,24,78,0,0,0,
102,78,0,110,106,0,109,0,99,25,64,0,0,0,
66,55,86,48,0,81,0,57,58,91,0,68,0,0,
45,8,37,0,105,74,30,111,0,52,0,84,0,0,
51,51,106,0,54,37,82,0,107,0,85,26,0,0,
77,108,118,25,19,0,72,0,62,17,0,0,0,0,
100,19,36,76,66,0,0,59,99,4,0,32,0,0,
0,18,69,49,55,88,0,58,101,0,63,26,0,0,
77,108,119,25,19,0,72,0,62,18,1,0,0,0,
26,97,101,62,85,0,10,17,0,37,0,82,0,0,
13,0,67,4,56,106,110,26,0,0,113,57,0,0,
13,0,68,4,56,106,111,27,0,0,113,57,0,0,
20,65,2,0,102,112,89,36,0,23,77,0,0,0,
0,74,91,17,116,23,33,0,69,0,65,99,0,0,
109,76,95,65,91,0,16,79,0,18,0,73,0,0,
106,74,64,39,69,0,60,0,85,10,88,0,0,0,
108,94,0,46,11,88,0,107,63,63,0,72,0,0,
12,8,88,89,0,101,110,27,0,43,0,13,0,0,
102,78,119,109,105,0,109,0,99,25,63,0,0,0,
0,93,117,105,14,60,0,31,50,0,10,60,0,0,
81,66,62,0,53,112,6,58,0,91,28,0,0,0,
0,73,90,17,116,23,0,32,68,0,65,98,0,0,
32,48,2,22,0,100,1,0,109,0,75,56,0,0,
21,95,11,0,12,49,0,55,5,0,23,38,0,0,
0,27,70,60,67,15,100,0,91,0,54,21,0,0,
96,61,84,0,101,17,9,0,49,95,0,62,0,0,
44,43,52,40,13,0,16,47,0,0,17,35,0,0,
74,84,34,16,0,19,0,6,98,63,0,25,0,0,
82,66,62,54,0,112,6,58,0,91,28,0,0,0,
17,72,40,90,0,25,0,116,111,0,29,90,0,0,
96,61,84,0,101,17,8,0,49,94,0,62,0,0,
21,95,11,0,13,49,0,56,5,0,23,38,0,0,
45,9,38,0,105,74,31,111,0,52,0,85,0,0,
0,73,91,17,116,23,33,0,68,0,65,99,0,0,
66,54,85,47,0,81,0,57,57,91,0,67,0,0,
67,56,4,68,0,57,89,0,23,58,0,17,0,0,
12,7,87,89,0,100,109,26,0,43,0,12,0,0,
17,113,38,0,64,75,46,0,85,0,107,13,0,0,
114,80,78,0,32,64,108,0,28,101,0,30,0,0,
7,84,71,0,93,116,0,60,5,32,107,0,0,0,
51,58,62,115,0,34,30,38,0,77,0,61,0,0,
0,26,70,60,67,15,100,0,91,0,54,20,0,0,
44,44,53,40,13,0,16,48,0,0,18,35,0,0,
118,114,55,15,98,0,26,53,0,60,84,0,0,0,
33,48,2,22,0,100,1,0,110,0,75,57,0,0,
111,31,71,0,13,74,0,76,6,93,0,101,0,0,
		others => 0);
	end function;
end package body;
